//////////////////////////////////////////////////////////////////////////////////////////
// Authors:      Alessandra Dolmeta - alessandra.dolmeta@polito.it                      //
//               Valeria Piscopo    - valeria.piscopo@polito.it                         //
//               Mattia Mirigaldi    - mattia.mirigaldi@polito.it                       //
// Language:     SystemVerilog                                                          //
// Based on the designed of Michal Peeters and Gilles Van Assche.                       //
//                                                                                      //
//////////////////////////////////////////////////////////////////////////////////////////

// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package keccak_reg_pkg;

  // Address widths within the block
  parameter int BlockAw = 8;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    logic [31:0] q;
  } keccak_reg2hw_data_mreg_t;

  typedef struct packed {
    logic        q;
  } keccak_reg2hw_ctrl_reg_t;

  typedef struct packed {
    logic [31:0] d;
    logic        de;
  } keccak_hw2reg_data_mreg_t;

  typedef struct packed {
    logic        d;
    logic        de;
  } keccak_hw2reg_status_reg_t;

  // Register -> HW type
  typedef struct packed {
    keccak_reg2hw_data_mreg_t [49:0] data; // [1600:1]
    keccak_reg2hw_ctrl_reg_t ctrl; // [0:0]
  } keccak_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    keccak_hw2reg_data_mreg_t [49:0] data; // [1651:2]
    keccak_hw2reg_status_reg_t status; // [1:0]
  } keccak_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] KECCAK_DATA_0_OFFSET = 8'h 0;
  parameter logic [BlockAw-1:0] KECCAK_DATA_1_OFFSET = 8'h 4;
  parameter logic [BlockAw-1:0] KECCAK_DATA_2_OFFSET = 8'h 8;
  parameter logic [BlockAw-1:0] KECCAK_DATA_3_OFFSET = 8'h c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_4_OFFSET = 8'h 10;
  parameter logic [BlockAw-1:0] KECCAK_DATA_5_OFFSET = 8'h 14;
  parameter logic [BlockAw-1:0] KECCAK_DATA_6_OFFSET = 8'h 18;
  parameter logic [BlockAw-1:0] KECCAK_DATA_7_OFFSET = 8'h 1c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_8_OFFSET = 8'h 20;
  parameter logic [BlockAw-1:0] KECCAK_DATA_9_OFFSET = 8'h 24;
  parameter logic [BlockAw-1:0] KECCAK_DATA_10_OFFSET = 8'h 28;
  parameter logic [BlockAw-1:0] KECCAK_DATA_11_OFFSET = 8'h 2c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_12_OFFSET = 8'h 30;
  parameter logic [BlockAw-1:0] KECCAK_DATA_13_OFFSET = 8'h 34;
  parameter logic [BlockAw-1:0] KECCAK_DATA_14_OFFSET = 8'h 38;
  parameter logic [BlockAw-1:0] KECCAK_DATA_15_OFFSET = 8'h 3c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_16_OFFSET = 8'h 40;
  parameter logic [BlockAw-1:0] KECCAK_DATA_17_OFFSET = 8'h 44;
  parameter logic [BlockAw-1:0] KECCAK_DATA_18_OFFSET = 8'h 48;
  parameter logic [BlockAw-1:0] KECCAK_DATA_19_OFFSET = 8'h 4c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_20_OFFSET = 8'h 50;
  parameter logic [BlockAw-1:0] KECCAK_DATA_21_OFFSET = 8'h 54;
  parameter logic [BlockAw-1:0] KECCAK_DATA_22_OFFSET = 8'h 58;
  parameter logic [BlockAw-1:0] KECCAK_DATA_23_OFFSET = 8'h 5c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_24_OFFSET = 8'h 60;
  parameter logic [BlockAw-1:0] KECCAK_DATA_25_OFFSET = 8'h 64;
  parameter logic [BlockAw-1:0] KECCAK_DATA_26_OFFSET = 8'h 68;
  parameter logic [BlockAw-1:0] KECCAK_DATA_27_OFFSET = 8'h 6c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_28_OFFSET = 8'h 70;
  parameter logic [BlockAw-1:0] KECCAK_DATA_29_OFFSET = 8'h 74;
  parameter logic [BlockAw-1:0] KECCAK_DATA_30_OFFSET = 8'h 78;
  parameter logic [BlockAw-1:0] KECCAK_DATA_31_OFFSET = 8'h 7c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_32_OFFSET = 8'h 80;
  parameter logic [BlockAw-1:0] KECCAK_DATA_33_OFFSET = 8'h 84;
  parameter logic [BlockAw-1:0] KECCAK_DATA_34_OFFSET = 8'h 88;
  parameter logic [BlockAw-1:0] KECCAK_DATA_35_OFFSET = 8'h 8c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_36_OFFSET = 8'h 90;
  parameter logic [BlockAw-1:0] KECCAK_DATA_37_OFFSET = 8'h 94;
  parameter logic [BlockAw-1:0] KECCAK_DATA_38_OFFSET = 8'h 98;
  parameter logic [BlockAw-1:0] KECCAK_DATA_39_OFFSET = 8'h 9c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_40_OFFSET = 8'h a0;
  parameter logic [BlockAw-1:0] KECCAK_DATA_41_OFFSET = 8'h a4;
  parameter logic [BlockAw-1:0] KECCAK_DATA_42_OFFSET = 8'h a8;
  parameter logic [BlockAw-1:0] KECCAK_DATA_43_OFFSET = 8'h ac;
  parameter logic [BlockAw-1:0] KECCAK_DATA_44_OFFSET = 8'h b0;
  parameter logic [BlockAw-1:0] KECCAK_DATA_45_OFFSET = 8'h b4;
  parameter logic [BlockAw-1:0] KECCAK_DATA_46_OFFSET = 8'h b8;
  parameter logic [BlockAw-1:0] KECCAK_DATA_47_OFFSET = 8'h bc;
  parameter logic [BlockAw-1:0] KECCAK_DATA_48_OFFSET = 8'h c0;
  parameter logic [BlockAw-1:0] KECCAK_DATA_49_OFFSET = 8'h c4;
  parameter logic [BlockAw-1:0] KECCAK_CTRL_OFFSET = 8'h c8;
  parameter logic [BlockAw-1:0] KECCAK_STATUS_OFFSET = 8'h cc;

  // Register index
  typedef enum int {
    KECCAK_DATA_0,
    KECCAK_DATA_1,
    KECCAK_DATA_2,
    KECCAK_DATA_3,
    KECCAK_DATA_4,
    KECCAK_DATA_5,
    KECCAK_DATA_6,
    KECCAK_DATA_7,
    KECCAK_DATA_8,
    KECCAK_DATA_9,
    KECCAK_DATA_10,
    KECCAK_DATA_11,
    KECCAK_DATA_12,
    KECCAK_DATA_13,
    KECCAK_DATA_14,
    KECCAK_DATA_15,
    KECCAK_DATA_16,
    KECCAK_DATA_17,
    KECCAK_DATA_18,
    KECCAK_DATA_19,
    KECCAK_DATA_20,
    KECCAK_DATA_21,
    KECCAK_DATA_22,
    KECCAK_DATA_23,
    KECCAK_DATA_24,
    KECCAK_DATA_25,
    KECCAK_DATA_26,
    KECCAK_DATA_27,
    KECCAK_DATA_28,
    KECCAK_DATA_29,
    KECCAK_DATA_30,
    KECCAK_DATA_31,
    KECCAK_DATA_32,
    KECCAK_DATA_33,
    KECCAK_DATA_34,
    KECCAK_DATA_35,
    KECCAK_DATA_36,
    KECCAK_DATA_37,
    KECCAK_DATA_38,
    KECCAK_DATA_39,
    KECCAK_DATA_40,
    KECCAK_DATA_41,
    KECCAK_DATA_42,
    KECCAK_DATA_43,
    KECCAK_DATA_44,
    KECCAK_DATA_45,
    KECCAK_DATA_46,
    KECCAK_DATA_47,
    KECCAK_DATA_48,
    KECCAK_DATA_49,
    KECCAK_CTRL,
    KECCAK_STATUS
  } keccak_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] KECCAK_PERMIT [52] = '{
    4'b 1111, // index[ 0] KECCAK_DATA_0
    4'b 1111, // index[ 1] KECCAK_DATA_1
    4'b 1111, // index[ 2] KECCAK_DATA_2
    4'b 1111, // index[ 3] KECCAK_DATA_3
    4'b 1111, // index[ 4] KECCAK_DATA_4
    4'b 1111, // index[ 5] KECCAK_DATA_5
    4'b 1111, // index[ 6] KECCAK_DATA_6
    4'b 1111, // index[ 7] KECCAK_DATA_7
    4'b 1111, // index[ 8] KECCAK_DATA_8
    4'b 1111, // index[ 9] KECCAK_DATA_9
    4'b 1111, // index[10] KECCAK_DATA_10
    4'b 1111, // index[11] KECCAK_DATA_11
    4'b 1111, // index[12] KECCAK_DATA_12
    4'b 1111, // index[13] KECCAK_DATA_13
    4'b 1111, // index[14] KECCAK_DATA_14
    4'b 1111, // index[15] KECCAK_DATA_15
    4'b 1111, // index[16] KECCAK_DATA_16
    4'b 1111, // index[17] KECCAK_DATA_17
    4'b 1111, // index[18] KECCAK_DATA_18
    4'b 1111, // index[19] KECCAK_DATA_19
    4'b 1111, // index[20] KECCAK_DATA_20
    4'b 1111, // index[21] KECCAK_DATA_21
    4'b 1111, // index[22] KECCAK_DATA_22
    4'b 1111, // index[23] KECCAK_DATA_23
    4'b 1111, // index[24] KECCAK_DATA_24
    4'b 1111, // index[25] KECCAK_DATA_25
    4'b 1111, // index[26] KECCAK_DATA_26
    4'b 1111, // index[27] KECCAK_DATA_27
    4'b 1111, // index[28] KECCAK_DATA_28
    4'b 1111, // index[29] KECCAK_DATA_29
    4'b 1111, // index[30] KECCAK_DATA_30
    4'b 1111, // index[31] KECCAK_DATA_31
    4'b 1111, // index[32] KECCAK_DATA_32
    4'b 1111, // index[33] KECCAK_DATA_33
    4'b 1111, // index[34] KECCAK_DATA_34
    4'b 1111, // index[35] KECCAK_DATA_35
    4'b 1111, // index[36] KECCAK_DATA_36
    4'b 1111, // index[37] KECCAK_DATA_37
    4'b 1111, // index[38] KECCAK_DATA_38
    4'b 1111, // index[39] KECCAK_DATA_39
    4'b 1111, // index[40] KECCAK_DATA_40
    4'b 1111, // index[41] KECCAK_DATA_41
    4'b 1111, // index[42] KECCAK_DATA_42
    4'b 1111, // index[43] KECCAK_DATA_43
    4'b 1111, // index[44] KECCAK_DATA_44
    4'b 1111, // index[45] KECCAK_DATA_45
    4'b 1111, // index[46] KECCAK_DATA_46
    4'b 1111, // index[47] KECCAK_DATA_47
    4'b 1111, // index[48] KECCAK_DATA_48
    4'b 1111, // index[49] KECCAK_DATA_49
    4'b 0001, // index[50] KECCAK_CTRL
    4'b 0001  // index[51] KECCAK_STATUS
  };

endpackage

