//////////////////////////////////////////////////////////////////////////////////////////
// Authors:      Alessandra Dolmeta - alessandra.dolmeta@polito.it                      //
//               Valeria Piscopo    - valeria.piscopo@polito.it                         //
//               Mattia Mirigaldi    - mattia.mirigaldi@polito.it                       //
// Language:     SystemVerilog                                                          //
// Based on the designed of Michal Peeters and Gilles Van Assche.                       //
//                                                                                      //
//////////////////////////////////////////////////////////////////////////////////////////

// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`


`include "common_cells/assertions.svh"

module keccak_reg_top #(
  parameter type reg_req_t = logic,
  parameter type reg_rsp_t = logic,
  parameter int AW = 8
) (
  input logic clk_i,
  input logic rst_ni,
  input  reg_req_t reg_req_i,
  output reg_rsp_t reg_rsp_o,
  // To HW
  output keccak_reg_pkg::keccak_reg2hw_t reg2hw, // Write
  input  keccak_reg_pkg::keccak_hw2reg_t hw2reg, // Read


  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import keccak_reg_pkg::* ;

  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;

  // Below register interface can be changed
  reg_req_t  reg_intf_req;
  reg_rsp_t  reg_intf_rsp;


  assign reg_intf_req = reg_req_i;
  assign reg_rsp_o = reg_intf_rsp;


  assign reg_we = reg_intf_req.valid & reg_intf_req.write;
  assign reg_re = reg_intf_req.valid & ~reg_intf_req.write;
  assign reg_addr = reg_intf_req.addr;
  assign reg_wdata = reg_intf_req.wdata;
  assign reg_be = reg_intf_req.wstrb;
  assign reg_intf_rsp.rdata = reg_rdata;
  assign reg_intf_rsp.error = reg_error;
  assign reg_intf_rsp.ready = 1'b1;

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err;


  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic [31:0] data_0_qs;
  logic [31:0] data_0_wd;
  logic data_0_we;
  logic [31:0] data_1_qs;
  logic [31:0] data_1_wd;
  logic data_1_we;
  logic [31:0] data_2_qs;
  logic [31:0] data_2_wd;
  logic data_2_we;
  logic [31:0] data_3_qs;
  logic [31:0] data_3_wd;
  logic data_3_we;
  logic [31:0] data_4_qs;
  logic [31:0] data_4_wd;
  logic data_4_we;
  logic [31:0] data_5_qs;
  logic [31:0] data_5_wd;
  logic data_5_we;
  logic [31:0] data_6_qs;
  logic [31:0] data_6_wd;
  logic data_6_we;
  logic [31:0] data_7_qs;
  logic [31:0] data_7_wd;
  logic data_7_we;
  logic [31:0] data_8_qs;
  logic [31:0] data_8_wd;
  logic data_8_we;
  logic [31:0] data_9_qs;
  logic [31:0] data_9_wd;
  logic data_9_we;
  logic [31:0] data_10_qs;
  logic [31:0] data_10_wd;
  logic data_10_we;
  logic [31:0] data_11_qs;
  logic [31:0] data_11_wd;
  logic data_11_we;
  logic [31:0] data_12_qs;
  logic [31:0] data_12_wd;
  logic data_12_we;
  logic [31:0] data_13_qs;
  logic [31:0] data_13_wd;
  logic data_13_we;
  logic [31:0] data_14_qs;
  logic [31:0] data_14_wd;
  logic data_14_we;
  logic [31:0] data_15_qs;
  logic [31:0] data_15_wd;
  logic data_15_we;
  logic [31:0] data_16_qs;
  logic [31:0] data_16_wd;
  logic data_16_we;
  logic [31:0] data_17_qs;
  logic [31:0] data_17_wd;
  logic data_17_we;
  logic [31:0] data_18_qs;
  logic [31:0] data_18_wd;
  logic data_18_we;
  logic [31:0] data_19_qs;
  logic [31:0] data_19_wd;
  logic data_19_we;
  logic [31:0] data_20_qs;
  logic [31:0] data_20_wd;
  logic data_20_we;
  logic [31:0] data_21_qs;
  logic [31:0] data_21_wd;
  logic data_21_we;
  logic [31:0] data_22_qs;
  logic [31:0] data_22_wd;
  logic data_22_we;
  logic [31:0] data_23_qs;
  logic [31:0] data_23_wd;
  logic data_23_we;
  logic [31:0] data_24_qs;
  logic [31:0] data_24_wd;
  logic data_24_we;
  logic [31:0] data_25_qs;
  logic [31:0] data_25_wd;
  logic data_25_we;
  logic [31:0] data_26_qs;
  logic [31:0] data_26_wd;
  logic data_26_we;
  logic [31:0] data_27_qs;
  logic [31:0] data_27_wd;
  logic data_27_we;
  logic [31:0] data_28_qs;
  logic [31:0] data_28_wd;
  logic data_28_we;
  logic [31:0] data_29_qs;
  logic [31:0] data_29_wd;
  logic data_29_we;
  logic [31:0] data_30_qs;
  logic [31:0] data_30_wd;
  logic data_30_we;
  logic [31:0] data_31_qs;
  logic [31:0] data_31_wd;
  logic data_31_we;
  logic [31:0] data_32_qs;
  logic [31:0] data_32_wd;
  logic data_32_we;
  logic [31:0] data_33_qs;
  logic [31:0] data_33_wd;
  logic data_33_we;
  logic [31:0] data_34_qs;
  logic [31:0] data_34_wd;
  logic data_34_we;
  logic [31:0] data_35_qs;
  logic [31:0] data_35_wd;
  logic data_35_we;
  logic [31:0] data_36_qs;
  logic [31:0] data_36_wd;
  logic data_36_we;
  logic [31:0] data_37_qs;
  logic [31:0] data_37_wd;
  logic data_37_we;
  logic [31:0] data_38_qs;
  logic [31:0] data_38_wd;
  logic data_38_we;
  logic [31:0] data_39_qs;
  logic [31:0] data_39_wd;
  logic data_39_we;
  logic [31:0] data_40_qs;
  logic [31:0] data_40_wd;
  logic data_40_we;
  logic [31:0] data_41_qs;
  logic [31:0] data_41_wd;
  logic data_41_we;
  logic [31:0] data_42_qs;
  logic [31:0] data_42_wd;
  logic data_42_we;
  logic [31:0] data_43_qs;
  logic [31:0] data_43_wd;
  logic data_43_we;
  logic [31:0] data_44_qs;
  logic [31:0] data_44_wd;
  logic data_44_we;
  logic [31:0] data_45_qs;
  logic [31:0] data_45_wd;
  logic data_45_we;
  logic [31:0] data_46_qs;
  logic [31:0] data_46_wd;
  logic data_46_we;
  logic [31:0] data_47_qs;
  logic [31:0] data_47_wd;
  logic data_47_we;
  logic [31:0] data_48_qs;
  logic [31:0] data_48_wd;
  logic data_48_we;
  logic [31:0] data_49_qs;
  logic [31:0] data_49_wd;
  logic data_49_we;
  logic ctrl_wd;
  logic ctrl_we;
  logic status_qs;

  // Register instances

  // Subregister 0 of Multireg data
  // R[data_0]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_0 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_0_we),
    .wd     (data_0_wd),

    // from internal hardware
    .de     (hw2reg.data[0].de),
    .d      (hw2reg.data[0].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[0].q ),

    // to register interface (read)
    .qs     (data_0_qs)
  );

  // Subregister 1 of Multireg data
  // R[data_1]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_1 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_1_we),
    .wd     (data_1_wd),

    // from internal hardware
    .de     (hw2reg.data[1].de),
    .d      (hw2reg.data[1].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[1].q ),

    // to register interface (read)
    .qs     (data_1_qs)
  );

  // Subregister 2 of Multireg data
  // R[data_2]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_2 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_2_we),
    .wd     (data_2_wd),

    // from internal hardware
    .de     (hw2reg.data[2].de),
    .d      (hw2reg.data[2].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[2].q ),

    // to register interface (read)
    .qs     (data_2_qs)
  );

  // Subregister 3 of Multireg data
  // R[data_3]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_3 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_3_we),
    .wd     (data_3_wd),

    // from internal hardware
    .de     (hw2reg.data[3].de),
    .d      (hw2reg.data[3].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[3].q ),

    // to register interface (read)
    .qs     (data_3_qs)
  );

  // Subregister 4 of Multireg data
  // R[data_4]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_4 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_4_we),
    .wd     (data_4_wd),

    // from internal hardware
    .de     (hw2reg.data[4].de),
    .d      (hw2reg.data[4].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[4].q ),

    // to register interface (read)
    .qs     (data_4_qs)
  );

  // Subregister 5 of Multireg data
  // R[data_5]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_5 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_5_we),
    .wd     (data_5_wd),

    // from internal hardware
    .de     (hw2reg.data[5].de),
    .d      (hw2reg.data[5].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[5].q ),

    // to register interface (read)
    .qs     (data_5_qs)
  );

  // Subregister 6 of Multireg data
  // R[data_6]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_6 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_6_we),
    .wd     (data_6_wd),

    // from internal hardware
    .de     (hw2reg.data[6].de),
    .d      (hw2reg.data[6].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[6].q ),

    // to register interface (read)
    .qs     (data_6_qs)
  );

  // Subregister 7 of Multireg data
  // R[data_7]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_7 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_7_we),
    .wd     (data_7_wd),

    // from internal hardware
    .de     (hw2reg.data[7].de),
    .d      (hw2reg.data[7].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[7].q ),

    // to register interface (read)
    .qs     (data_7_qs)
  );

  // Subregister 8 of Multireg data
  // R[data_8]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_8 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_8_we),
    .wd     (data_8_wd),

    // from internal hardware
    .de     (hw2reg.data[8].de),
    .d      (hw2reg.data[8].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[8].q ),

    // to register interface (read)
    .qs     (data_8_qs)
  );

  // Subregister 9 of Multireg data
  // R[data_9]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_9 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_9_we),
    .wd     (data_9_wd),

    // from internal hardware
    .de     (hw2reg.data[9].de),
    .d      (hw2reg.data[9].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[9].q ),

    // to register interface (read)
    .qs     (data_9_qs)
  );

  // Subregister 10 of Multireg data
  // R[data_10]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_10 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_10_we),
    .wd     (data_10_wd),

    // from internal hardware
    .de     (hw2reg.data[10].de),
    .d      (hw2reg.data[10].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[10].q ),

    // to register interface (read)
    .qs     (data_10_qs)
  );

  // Subregister 11 of Multireg data
  // R[data_11]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_11 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_11_we),
    .wd     (data_11_wd),

    // from internal hardware
    .de     (hw2reg.data[11].de),
    .d      (hw2reg.data[11].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[11].q ),

    // to register interface (read)
    .qs     (data_11_qs)
  );

  // Subregister 12 of Multireg data
  // R[data_12]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_12 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_12_we),
    .wd     (data_12_wd),

    // from internal hardware
    .de     (hw2reg.data[12].de),
    .d      (hw2reg.data[12].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[12].q ),

    // to register interface (read)
    .qs     (data_12_qs)
  );

  // Subregister 13 of Multireg data
  // R[data_13]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_13 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_13_we),
    .wd     (data_13_wd),

    // from internal hardware
    .de     (hw2reg.data[13].de),
    .d      (hw2reg.data[13].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[13].q ),

    // to register interface (read)
    .qs     (data_13_qs)
  );

  // Subregister 14 of Multireg data
  // R[data_14]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_14 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_14_we),
    .wd     (data_14_wd),

    // from internal hardware
    .de     (hw2reg.data[14].de),
    .d      (hw2reg.data[14].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[14].q ),

    // to register interface (read)
    .qs     (data_14_qs)
  );

  // Subregister 15 of Multireg data
  // R[data_15]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_15 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_15_we),
    .wd     (data_15_wd),

    // from internal hardware
    .de     (hw2reg.data[15].de),
    .d      (hw2reg.data[15].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[15].q ),

    // to register interface (read)
    .qs     (data_15_qs)
  );

  // Subregister 16 of Multireg data
  // R[data_16]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_16 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_16_we),
    .wd     (data_16_wd),

    // from internal hardware
    .de     (hw2reg.data[16].de),
    .d      (hw2reg.data[16].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[16].q ),

    // to register interface (read)
    .qs     (data_16_qs)
  );

  // Subregister 17 of Multireg data
  // R[data_17]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_17 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_17_we),
    .wd     (data_17_wd),

    // from internal hardware
    .de     (hw2reg.data[17].de),
    .d      (hw2reg.data[17].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[17].q ),

    // to register interface (read)
    .qs     (data_17_qs)
  );

  // Subregister 18 of Multireg data
  // R[data_18]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_18 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_18_we),
    .wd     (data_18_wd),

    // from internal hardware
    .de     (hw2reg.data[18].de),
    .d      (hw2reg.data[18].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[18].q ),

    // to register interface (read)
    .qs     (data_18_qs)
  );

  // Subregister 19 of Multireg data
  // R[data_19]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_19 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_19_we),
    .wd     (data_19_wd),

    // from internal hardware
    .de     (hw2reg.data[19].de),
    .d      (hw2reg.data[19].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[19].q ),

    // to register interface (read)
    .qs     (data_19_qs)
  );

  // Subregister 20 of Multireg data
  // R[data_20]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_20 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_20_we),
    .wd     (data_20_wd),

    // from internal hardware
    .de     (hw2reg.data[20].de),
    .d      (hw2reg.data[20].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[20].q ),

    // to register interface (read)
    .qs     (data_20_qs)
  );

  // Subregister 21 of Multireg data
  // R[data_21]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_21 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_21_we),
    .wd     (data_21_wd),

    // from internal hardware
    .de     (hw2reg.data[21].de),
    .d      (hw2reg.data[21].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[21].q ),

    // to register interface (read)
    .qs     (data_21_qs)
  );

  // Subregister 22 of Multireg data
  // R[data_22]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_22 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_22_we),
    .wd     (data_22_wd),

    // from internal hardware
    .de     (hw2reg.data[22].de),
    .d      (hw2reg.data[22].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[22].q ),

    // to register interface (read)
    .qs     (data_22_qs)
  );

  // Subregister 23 of Multireg data
  // R[data_23]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_23 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_23_we),
    .wd     (data_23_wd),

    // from internal hardware
    .de     (hw2reg.data[23].de),
    .d      (hw2reg.data[23].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[23].q ),

    // to register interface (read)
    .qs     (data_23_qs)
  );

  // Subregister 24 of Multireg data
  // R[data_24]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_24 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_24_we),
    .wd     (data_24_wd),

    // from internal hardware
    .de     (hw2reg.data[24].de),
    .d      (hw2reg.data[24].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[24].q ),

    // to register interface (read)
    .qs     (data_24_qs)
  );

  // Subregister 25 of Multireg data
  // R[data_25]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_25 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_25_we),
    .wd     (data_25_wd),

    // from internal hardware
    .de     (hw2reg.data[25].de),
    .d      (hw2reg.data[25].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[25].q ),

    // to register interface (read)
    .qs     (data_25_qs)
  );

  // Subregister 26 of Multireg data
  // R[data_26]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_26 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_26_we),
    .wd     (data_26_wd),

    // from internal hardware
    .de     (hw2reg.data[26].de),
    .d      (hw2reg.data[26].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[26].q ),

    // to register interface (read)
    .qs     (data_26_qs)
  );

  // Subregister 27 of Multireg data
  // R[data_27]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_27 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_27_we),
    .wd     (data_27_wd),

    // from internal hardware
    .de     (hw2reg.data[27].de),
    .d      (hw2reg.data[27].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[27].q ),

    // to register interface (read)
    .qs     (data_27_qs)
  );

  // Subregister 28 of Multireg data
  // R[data_28]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_28 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_28_we),
    .wd     (data_28_wd),

    // from internal hardware
    .de     (hw2reg.data[28].de),
    .d      (hw2reg.data[28].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[28].q ),

    // to register interface (read)
    .qs     (data_28_qs)
  );

  // Subregister 29 of Multireg data
  // R[data_29]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_29 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_29_we),
    .wd     (data_29_wd),

    // from internal hardware
    .de     (hw2reg.data[29].de),
    .d      (hw2reg.data[29].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[29].q ),

    // to register interface (read)
    .qs     (data_29_qs)
  );

  // Subregister 30 of Multireg data
  // R[data_30]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_30 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_30_we),
    .wd     (data_30_wd),

    // from internal hardware
    .de     (hw2reg.data[30].de),
    .d      (hw2reg.data[30].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[30].q ),

    // to register interface (read)
    .qs     (data_30_qs)
  );

  // Subregister 31 of Multireg data
  // R[data_31]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_31 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_31_we),
    .wd     (data_31_wd),

    // from internal hardware
    .de     (hw2reg.data[31].de),
    .d      (hw2reg.data[31].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[31].q ),

    // to register interface (read)
    .qs     (data_31_qs)
  );

  // Subregister 32 of Multireg data
  // R[data_32]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_32 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_32_we),
    .wd     (data_32_wd),

    // from internal hardware
    .de     (hw2reg.data[32].de),
    .d      (hw2reg.data[32].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[32].q ),

    // to register interface (read)
    .qs     (data_32_qs)
  );

  // Subregister 33 of Multireg data
  // R[data_33]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_33 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_33_we),
    .wd     (data_33_wd),

    // from internal hardware
    .de     (hw2reg.data[33].de),
    .d      (hw2reg.data[33].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[33].q ),

    // to register interface (read)
    .qs     (data_33_qs)
  );

  // Subregister 34 of Multireg data
  // R[data_34]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_34 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_34_we),
    .wd     (data_34_wd),

    // from internal hardware
    .de     (hw2reg.data[34].de),
    .d      (hw2reg.data[34].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[34].q ),

    // to register interface (read)
    .qs     (data_34_qs)
  );

  // Subregister 35 of Multireg data
  // R[data_35]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_35 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_35_we),
    .wd     (data_35_wd),

    // from internal hardware
    .de     (hw2reg.data[35].de),
    .d      (hw2reg.data[35].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[35].q ),

    // to register interface (read)
    .qs     (data_35_qs)
  );

  // Subregister 36 of Multireg data
  // R[data_36]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_36 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_36_we),
    .wd     (data_36_wd),

    // from internal hardware
    .de     (hw2reg.data[36].de),
    .d      (hw2reg.data[36].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[36].q ),

    // to register interface (read)
    .qs     (data_36_qs)
  );

  // Subregister 37 of Multireg data
  // R[data_37]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_37 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_37_we),
    .wd     (data_37_wd),

    // from internal hardware
    .de     (hw2reg.data[37].de),
    .d      (hw2reg.data[37].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[37].q ),

    // to register interface (read)
    .qs     (data_37_qs)
  );

  // Subregister 38 of Multireg data
  // R[data_38]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_38 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_38_we),
    .wd     (data_38_wd),

    // from internal hardware
    .de     (hw2reg.data[38].de),
    .d      (hw2reg.data[38].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[38].q ),

    // to register interface (read)
    .qs     (data_38_qs)
  );

  // Subregister 39 of Multireg data
  // R[data_39]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_39 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_39_we),
    .wd     (data_39_wd),

    // from internal hardware
    .de     (hw2reg.data[39].de),
    .d      (hw2reg.data[39].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[39].q ),

    // to register interface (read)
    .qs     (data_39_qs)
  );

  // Subregister 40 of Multireg data
  // R[data_40]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_40 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_40_we),
    .wd     (data_40_wd),

    // from internal hardware
    .de     (hw2reg.data[40].de),
    .d      (hw2reg.data[40].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[40].q ),

    // to register interface (read)
    .qs     (data_40_qs)
  );

  // Subregister 41 of Multireg data
  // R[data_41]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_41 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_41_we),
    .wd     (data_41_wd),

    // from internal hardware
    .de     (hw2reg.data[41].de),
    .d      (hw2reg.data[41].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[41].q ),

    // to register interface (read)
    .qs     (data_41_qs)
  );

  // Subregister 42 of Multireg data
  // R[data_42]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_42 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_42_we),
    .wd     (data_42_wd),

    // from internal hardware
    .de     (hw2reg.data[42].de),
    .d      (hw2reg.data[42].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[42].q ),

    // to register interface (read)
    .qs     (data_42_qs)
  );

  // Subregister 43 of Multireg data
  // R[data_43]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_43 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_43_we),
    .wd     (data_43_wd),

    // from internal hardware
    .de     (hw2reg.data[43].de),
    .d      (hw2reg.data[43].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[43].q ),

    // to register interface (read)
    .qs     (data_43_qs)
  );

  // Subregister 44 of Multireg data
  // R[data_44]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_44 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_44_we),
    .wd     (data_44_wd),

    // from internal hardware
    .de     (hw2reg.data[44].de),
    .d      (hw2reg.data[44].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[44].q ),

    // to register interface (read)
    .qs     (data_44_qs)
  );

  // Subregister 45 of Multireg data
  // R[data_45]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_45 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_45_we),
    .wd     (data_45_wd),

    // from internal hardware
    .de     (hw2reg.data[45].de),
    .d      (hw2reg.data[45].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[45].q ),

    // to register interface (read)
    .qs     (data_45_qs)
  );

  // Subregister 46 of Multireg data
  // R[data_46]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_46 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_46_we),
    .wd     (data_46_wd),

    // from internal hardware
    .de     (hw2reg.data[46].de),
    .d      (hw2reg.data[46].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[46].q ),

    // to register interface (read)
    .qs     (data_46_qs)
  );

  // Subregister 47 of Multireg data
  // R[data_47]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_47 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_47_we),
    .wd     (data_47_wd),

    // from internal hardware
    .de     (hw2reg.data[47].de),
    .d      (hw2reg.data[47].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[47].q ),

    // to register interface (read)
    .qs     (data_47_qs)
  );

  // Subregister 48 of Multireg data
  // R[data_48]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_48 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_48_we),
    .wd     (data_48_wd),

    // from internal hardware
    .de     (hw2reg.data[48].de),
    .d      (hw2reg.data[48].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[48].q ),

    // to register interface (read)
    .qs     (data_48_qs)
  );

  // Subregister 49 of Multireg data
  // R[data_49]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("RW"),
    .RESVAL  (32'h0)
  ) u_data_49 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (data_49_we),
    .wd     (data_49_wd),

    // from internal hardware
    .de     (hw2reg.data[49].de),
    .d      (hw2reg.data[49].d ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.data[49].q ),

    // to register interface (read)
    .qs     (data_49_qs)
  );


  // R[ctrl]: V(False)

  prim_subreg #(
    .DW      (1),
    .SWACCESS("WO"),
    .RESVAL  (1'h0)
  ) u_ctrl (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (ctrl_we),
    .wd     (ctrl_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.ctrl.q ),

    .qs     ()
  );


  // R[status]: V(False)

  prim_subreg #(
    .DW      (1),
    .SWACCESS("RO"),
    .RESVAL  (1'h0)
  ) u_status (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    .we     (1'b0),
    .wd     ('0  ),

    // from internal hardware
    .de     (hw2reg.status.de),
    .d      (hw2reg.status.d ),

    // to internal hardware
    .qe     (),
    .q      (),

    // to register interface (read)
    .qs     (status_qs)
  );




  logic [51:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == KECCAK_DATA_0_OFFSET);
    addr_hit[ 1] = (reg_addr == KECCAK_DATA_1_OFFSET);
    addr_hit[ 2] = (reg_addr == KECCAK_DATA_2_OFFSET);
    addr_hit[ 3] = (reg_addr == KECCAK_DATA_3_OFFSET);
    addr_hit[ 4] = (reg_addr == KECCAK_DATA_4_OFFSET);
    addr_hit[ 5] = (reg_addr == KECCAK_DATA_5_OFFSET);
    addr_hit[ 6] = (reg_addr == KECCAK_DATA_6_OFFSET);
    addr_hit[ 7] = (reg_addr == KECCAK_DATA_7_OFFSET);
    addr_hit[ 8] = (reg_addr == KECCAK_DATA_8_OFFSET);
    addr_hit[ 9] = (reg_addr == KECCAK_DATA_9_OFFSET);
    addr_hit[10] = (reg_addr == KECCAK_DATA_10_OFFSET);
    addr_hit[11] = (reg_addr == KECCAK_DATA_11_OFFSET);
    addr_hit[12] = (reg_addr == KECCAK_DATA_12_OFFSET);
    addr_hit[13] = (reg_addr == KECCAK_DATA_13_OFFSET);
    addr_hit[14] = (reg_addr == KECCAK_DATA_14_OFFSET);
    addr_hit[15] = (reg_addr == KECCAK_DATA_15_OFFSET);
    addr_hit[16] = (reg_addr == KECCAK_DATA_16_OFFSET);
    addr_hit[17] = (reg_addr == KECCAK_DATA_17_OFFSET);
    addr_hit[18] = (reg_addr == KECCAK_DATA_18_OFFSET);
    addr_hit[19] = (reg_addr == KECCAK_DATA_19_OFFSET);
    addr_hit[20] = (reg_addr == KECCAK_DATA_20_OFFSET);
    addr_hit[21] = (reg_addr == KECCAK_DATA_21_OFFSET);
    addr_hit[22] = (reg_addr == KECCAK_DATA_22_OFFSET);
    addr_hit[23] = (reg_addr == KECCAK_DATA_23_OFFSET);
    addr_hit[24] = (reg_addr == KECCAK_DATA_24_OFFSET);
    addr_hit[25] = (reg_addr == KECCAK_DATA_25_OFFSET);
    addr_hit[26] = (reg_addr == KECCAK_DATA_26_OFFSET);
    addr_hit[27] = (reg_addr == KECCAK_DATA_27_OFFSET);
    addr_hit[28] = (reg_addr == KECCAK_DATA_28_OFFSET);
    addr_hit[29] = (reg_addr == KECCAK_DATA_29_OFFSET);
    addr_hit[30] = (reg_addr == KECCAK_DATA_30_OFFSET);
    addr_hit[31] = (reg_addr == KECCAK_DATA_31_OFFSET);
    addr_hit[32] = (reg_addr == KECCAK_DATA_32_OFFSET);
    addr_hit[33] = (reg_addr == KECCAK_DATA_33_OFFSET);
    addr_hit[34] = (reg_addr == KECCAK_DATA_34_OFFSET);
    addr_hit[35] = (reg_addr == KECCAK_DATA_35_OFFSET);
    addr_hit[36] = (reg_addr == KECCAK_DATA_36_OFFSET);
    addr_hit[37] = (reg_addr == KECCAK_DATA_37_OFFSET);
    addr_hit[38] = (reg_addr == KECCAK_DATA_38_OFFSET);
    addr_hit[39] = (reg_addr == KECCAK_DATA_39_OFFSET);
    addr_hit[40] = (reg_addr == KECCAK_DATA_40_OFFSET);
    addr_hit[41] = (reg_addr == KECCAK_DATA_41_OFFSET);
    addr_hit[42] = (reg_addr == KECCAK_DATA_42_OFFSET);
    addr_hit[43] = (reg_addr == KECCAK_DATA_43_OFFSET);
    addr_hit[44] = (reg_addr == KECCAK_DATA_44_OFFSET);
    addr_hit[45] = (reg_addr == KECCAK_DATA_45_OFFSET);
    addr_hit[46] = (reg_addr == KECCAK_DATA_46_OFFSET);
    addr_hit[47] = (reg_addr == KECCAK_DATA_47_OFFSET);
    addr_hit[48] = (reg_addr == KECCAK_DATA_48_OFFSET);
    addr_hit[49] = (reg_addr == KECCAK_DATA_49_OFFSET);
    addr_hit[50] = (reg_addr == KECCAK_CTRL_OFFSET);
    addr_hit[51] = (reg_addr == KECCAK_STATUS_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(KECCAK_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(KECCAK_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(KECCAK_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(KECCAK_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(KECCAK_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(KECCAK_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(KECCAK_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(KECCAK_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(KECCAK_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(KECCAK_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(KECCAK_PERMIT[10] & ~reg_be))) |
               (addr_hit[11] & (|(KECCAK_PERMIT[11] & ~reg_be))) |
               (addr_hit[12] & (|(KECCAK_PERMIT[12] & ~reg_be))) |
               (addr_hit[13] & (|(KECCAK_PERMIT[13] & ~reg_be))) |
               (addr_hit[14] & (|(KECCAK_PERMIT[14] & ~reg_be))) |
               (addr_hit[15] & (|(KECCAK_PERMIT[15] & ~reg_be))) |
               (addr_hit[16] & (|(KECCAK_PERMIT[16] & ~reg_be))) |
               (addr_hit[17] & (|(KECCAK_PERMIT[17] & ~reg_be))) |
               (addr_hit[18] & (|(KECCAK_PERMIT[18] & ~reg_be))) |
               (addr_hit[19] & (|(KECCAK_PERMIT[19] & ~reg_be))) |
               (addr_hit[20] & (|(KECCAK_PERMIT[20] & ~reg_be))) |
               (addr_hit[21] & (|(KECCAK_PERMIT[21] & ~reg_be))) |
               (addr_hit[22] & (|(KECCAK_PERMIT[22] & ~reg_be))) |
               (addr_hit[23] & (|(KECCAK_PERMIT[23] & ~reg_be))) |
               (addr_hit[24] & (|(KECCAK_PERMIT[24] & ~reg_be))) |
               (addr_hit[25] & (|(KECCAK_PERMIT[25] & ~reg_be))) |
               (addr_hit[26] & (|(KECCAK_PERMIT[26] & ~reg_be))) |
               (addr_hit[27] & (|(KECCAK_PERMIT[27] & ~reg_be))) |
               (addr_hit[28] & (|(KECCAK_PERMIT[28] & ~reg_be))) |
               (addr_hit[29] & (|(KECCAK_PERMIT[29] & ~reg_be))) |
               (addr_hit[30] & (|(KECCAK_PERMIT[30] & ~reg_be))) |
               (addr_hit[31] & (|(KECCAK_PERMIT[31] & ~reg_be))) |
               (addr_hit[32] & (|(KECCAK_PERMIT[32] & ~reg_be))) |
               (addr_hit[33] & (|(KECCAK_PERMIT[33] & ~reg_be))) |
               (addr_hit[34] & (|(KECCAK_PERMIT[34] & ~reg_be))) |
               (addr_hit[35] & (|(KECCAK_PERMIT[35] & ~reg_be))) |
               (addr_hit[36] & (|(KECCAK_PERMIT[36] & ~reg_be))) |
               (addr_hit[37] & (|(KECCAK_PERMIT[37] & ~reg_be))) |
               (addr_hit[38] & (|(KECCAK_PERMIT[38] & ~reg_be))) |
               (addr_hit[39] & (|(KECCAK_PERMIT[39] & ~reg_be))) |
               (addr_hit[40] & (|(KECCAK_PERMIT[40] & ~reg_be))) |
               (addr_hit[41] & (|(KECCAK_PERMIT[41] & ~reg_be))) |
               (addr_hit[42] & (|(KECCAK_PERMIT[42] & ~reg_be))) |
               (addr_hit[43] & (|(KECCAK_PERMIT[43] & ~reg_be))) |
               (addr_hit[44] & (|(KECCAK_PERMIT[44] & ~reg_be))) |
               (addr_hit[45] & (|(KECCAK_PERMIT[45] & ~reg_be))) |
               (addr_hit[46] & (|(KECCAK_PERMIT[46] & ~reg_be))) |
               (addr_hit[47] & (|(KECCAK_PERMIT[47] & ~reg_be))) |
               (addr_hit[48] & (|(KECCAK_PERMIT[48] & ~reg_be))) |
               (addr_hit[49] & (|(KECCAK_PERMIT[49] & ~reg_be))) |
               (addr_hit[50] & (|(KECCAK_PERMIT[50] & ~reg_be))) |
               (addr_hit[51] & (|(KECCAK_PERMIT[51] & ~reg_be)))));
  end

  assign data_0_we = addr_hit[0] & reg_we & !reg_error;
  assign data_0_wd = reg_wdata[31:0];

  assign data_1_we = addr_hit[1] & reg_we & !reg_error;
  assign data_1_wd = reg_wdata[31:0];

  assign data_2_we = addr_hit[2] & reg_we & !reg_error;
  assign data_2_wd = reg_wdata[31:0];

  assign data_3_we = addr_hit[3] & reg_we & !reg_error;
  assign data_3_wd = reg_wdata[31:0];

  assign data_4_we = addr_hit[4] & reg_we & !reg_error;
  assign data_4_wd = reg_wdata[31:0];

  assign data_5_we = addr_hit[5] & reg_we & !reg_error;
  assign data_5_wd = reg_wdata[31:0];

  assign data_6_we = addr_hit[6] & reg_we & !reg_error;
  assign data_6_wd = reg_wdata[31:0];

  assign data_7_we = addr_hit[7] & reg_we & !reg_error;
  assign data_7_wd = reg_wdata[31:0];

  assign data_8_we = addr_hit[8] & reg_we & !reg_error;
  assign data_8_wd = reg_wdata[31:0];

  assign data_9_we = addr_hit[9] & reg_we & !reg_error;
  assign data_9_wd = reg_wdata[31:0];

  assign data_10_we = addr_hit[10] & reg_we & !reg_error;
  assign data_10_wd = reg_wdata[31:0];

  assign data_11_we = addr_hit[11] & reg_we & !reg_error;
  assign data_11_wd = reg_wdata[31:0];

  assign data_12_we = addr_hit[12] & reg_we & !reg_error;
  assign data_12_wd = reg_wdata[31:0];

  assign data_13_we = addr_hit[13] & reg_we & !reg_error;
  assign data_13_wd = reg_wdata[31:0];

  assign data_14_we = addr_hit[14] & reg_we & !reg_error;
  assign data_14_wd = reg_wdata[31:0];

  assign data_15_we = addr_hit[15] & reg_we & !reg_error;
  assign data_15_wd = reg_wdata[31:0];

  assign data_16_we = addr_hit[16] & reg_we & !reg_error;
  assign data_16_wd = reg_wdata[31:0];

  assign data_17_we = addr_hit[17] & reg_we & !reg_error;
  assign data_17_wd = reg_wdata[31:0];

  assign data_18_we = addr_hit[18] & reg_we & !reg_error;
  assign data_18_wd = reg_wdata[31:0];

  assign data_19_we = addr_hit[19] & reg_we & !reg_error;
  assign data_19_wd = reg_wdata[31:0];

  assign data_20_we = addr_hit[20] & reg_we & !reg_error;
  assign data_20_wd = reg_wdata[31:0];

  assign data_21_we = addr_hit[21] & reg_we & !reg_error;
  assign data_21_wd = reg_wdata[31:0];

  assign data_22_we = addr_hit[22] & reg_we & !reg_error;
  assign data_22_wd = reg_wdata[31:0];

  assign data_23_we = addr_hit[23] & reg_we & !reg_error;
  assign data_23_wd = reg_wdata[31:0];

  assign data_24_we = addr_hit[24] & reg_we & !reg_error;
  assign data_24_wd = reg_wdata[31:0];

  assign data_25_we = addr_hit[25] & reg_we & !reg_error;
  assign data_25_wd = reg_wdata[31:0];

  assign data_26_we = addr_hit[26] & reg_we & !reg_error;
  assign data_26_wd = reg_wdata[31:0];

  assign data_27_we = addr_hit[27] & reg_we & !reg_error;
  assign data_27_wd = reg_wdata[31:0];

  assign data_28_we = addr_hit[28] & reg_we & !reg_error;
  assign data_28_wd = reg_wdata[31:0];

  assign data_29_we = addr_hit[29] & reg_we & !reg_error;
  assign data_29_wd = reg_wdata[31:0];

  assign data_30_we = addr_hit[30] & reg_we & !reg_error;
  assign data_30_wd = reg_wdata[31:0];

  assign data_31_we = addr_hit[31] & reg_we & !reg_error;
  assign data_31_wd = reg_wdata[31:0];

  assign data_32_we = addr_hit[32] & reg_we & !reg_error;
  assign data_32_wd = reg_wdata[31:0];

  assign data_33_we = addr_hit[33] & reg_we & !reg_error;
  assign data_33_wd = reg_wdata[31:0];

  assign data_34_we = addr_hit[34] & reg_we & !reg_error;
  assign data_34_wd = reg_wdata[31:0];

  assign data_35_we = addr_hit[35] & reg_we & !reg_error;
  assign data_35_wd = reg_wdata[31:0];

  assign data_36_we = addr_hit[36] & reg_we & !reg_error;
  assign data_36_wd = reg_wdata[31:0];

  assign data_37_we = addr_hit[37] & reg_we & !reg_error;
  assign data_37_wd = reg_wdata[31:0];

  assign data_38_we = addr_hit[38] & reg_we & !reg_error;
  assign data_38_wd = reg_wdata[31:0];

  assign data_39_we = addr_hit[39] & reg_we & !reg_error;
  assign data_39_wd = reg_wdata[31:0];

  assign data_40_we = addr_hit[40] & reg_we & !reg_error;
  assign data_40_wd = reg_wdata[31:0];

  assign data_41_we = addr_hit[41] & reg_we & !reg_error;
  assign data_41_wd = reg_wdata[31:0];

  assign data_42_we = addr_hit[42] & reg_we & !reg_error;
  assign data_42_wd = reg_wdata[31:0];

  assign data_43_we = addr_hit[43] & reg_we & !reg_error;
  assign data_43_wd = reg_wdata[31:0];

  assign data_44_we = addr_hit[44] & reg_we & !reg_error;
  assign data_44_wd = reg_wdata[31:0];

  assign data_45_we = addr_hit[45] & reg_we & !reg_error;
  assign data_45_wd = reg_wdata[31:0];

  assign data_46_we = addr_hit[46] & reg_we & !reg_error;
  assign data_46_wd = reg_wdata[31:0];

  assign data_47_we = addr_hit[47] & reg_we & !reg_error;
  assign data_47_wd = reg_wdata[31:0];

  assign data_48_we = addr_hit[48] & reg_we & !reg_error;
  assign data_48_wd = reg_wdata[31:0];

  assign data_49_we = addr_hit[49] & reg_we & !reg_error;
  assign data_49_wd = reg_wdata[31:0];

  assign ctrl_we = addr_hit[50] & reg_we & !reg_error;
  assign ctrl_wd = reg_wdata[0];

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[31:0] = hw2reg.data[0].d;
      end

      addr_hit[1]: begin
        reg_rdata_next[31:0] = hw2reg.data[1].d;
      end

      addr_hit[2]: begin
        reg_rdata_next[31:0] = hw2reg.data[2].d;
      end

      addr_hit[3]: begin
        reg_rdata_next[31:0] = hw2reg.data[3].d;
      end

      addr_hit[4]: begin
        reg_rdata_next[31:0] = hw2reg.data[4].d;
      end

      addr_hit[5]: begin
        reg_rdata_next[31:0] = hw2reg.data[5].d;
      end

      addr_hit[6]: begin
        reg_rdata_next[31:0] = hw2reg.data[6].d;
      end

      addr_hit[7]: begin
        reg_rdata_next[31:0] = hw2reg.data[7].d;
      end

      addr_hit[8]: begin
        reg_rdata_next[31:0] = hw2reg.data[8].d;
      end

      addr_hit[9]: begin
        reg_rdata_next[31:0] = hw2reg.data[9].d;
      end

      addr_hit[10]: begin
        reg_rdata_next[31:0] = hw2reg.data[10].d;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = hw2reg.data[11].d;
      end

      addr_hit[12]: begin
        reg_rdata_next[31:0] = hw2reg.data[12].d;
      end

      addr_hit[13]: begin
        reg_rdata_next[31:0] = hw2reg.data[13].d;
      end

      addr_hit[14]: begin
        reg_rdata_next[31:0] = hw2reg.data[14].d;
      end

      addr_hit[15]: begin
        reg_rdata_next[31:0] = hw2reg.data[15].d;
      end

      addr_hit[16]: begin
        reg_rdata_next[31:0] = hw2reg.data[16].d;
      end

      addr_hit[17]: begin
        reg_rdata_next[31:0] = hw2reg.data[17].d;
      end

      addr_hit[18]: begin
        reg_rdata_next[31:0] = hw2reg.data[18].d;
      end

      addr_hit[19]: begin
        reg_rdata_next[31:0] = hw2reg.data[19].d;
      end

      addr_hit[20]: begin
        reg_rdata_next[31:0] = hw2reg.data[20].d;
      end

      addr_hit[21]: begin
        reg_rdata_next[31:0] = hw2reg.data[21].d;
      end

      addr_hit[22]: begin
        reg_rdata_next[31:0] = hw2reg.data[22].d;
      end

      addr_hit[23]: begin
        reg_rdata_next[31:0] = hw2reg.data[23].d;
      end

      addr_hit[24]: begin
        reg_rdata_next[31:0] = hw2reg.data[24].d;
      end

      addr_hit[25]: begin
        reg_rdata_next[31:0] = hw2reg.data[25].d;
      end

      addr_hit[26]: begin
        reg_rdata_next[31:0] = hw2reg.data[26].d;
      end

      addr_hit[27]: begin
        reg_rdata_next[31:0] = hw2reg.data[27].d;
      end

      addr_hit[28]: begin
        reg_rdata_next[31:0] = hw2reg.data[28].d;
      end

      addr_hit[29]: begin
        reg_rdata_next[31:0] = hw2reg.data[29].d;
      end

      addr_hit[30]: begin
        reg_rdata_next[31:0] = hw2reg.data[30].d;
      end

      addr_hit[31]: begin
        reg_rdata_next[31:0] = hw2reg.data[31].d;
      end

      addr_hit[32]: begin
        reg_rdata_next[31:0] = hw2reg.data[32].d;
      end

      addr_hit[33]: begin
        reg_rdata_next[31:0] = hw2reg.data[33].d;
      end

      addr_hit[34]: begin
        reg_rdata_next[31:0] = hw2reg.data[34].d;
      end

      addr_hit[35]: begin
        reg_rdata_next[31:0] = hw2reg.data[35].d;
      end

      addr_hit[36]: begin
        reg_rdata_next[31:0] = hw2reg.data[36].d;
      end

      addr_hit[37]: begin
        reg_rdata_next[31:0] = hw2reg.data[37].d;
      end

      addr_hit[38]: begin
        reg_rdata_next[31:0] = hw2reg.data[38].d;
      end

      addr_hit[39]: begin
        reg_rdata_next[31:0] = hw2reg.data[39].d;
      end

      addr_hit[40]: begin
        reg_rdata_next[31:0] = hw2reg.data[40].d;
      end

      addr_hit[41]: begin
        reg_rdata_next[31:0] = hw2reg.data[41].d;
      end

      addr_hit[42]: begin
        reg_rdata_next[31:0] = hw2reg.data[42].d;
      end

      addr_hit[43]: begin
        reg_rdata_next[31:0] = hw2reg.data[43].d;
      end

      addr_hit[44]: begin
        reg_rdata_next[31:0] = hw2reg.data[44].d;
      end

      addr_hit[45]: begin
        reg_rdata_next[31:0] = hw2reg.data[45].d;
      end

      addr_hit[46]: begin
        reg_rdata_next[31:0] = hw2reg.data[46].d;
      end

      addr_hit[47]: begin
        reg_rdata_next[31:0] = hw2reg.data[47].d;
      end

      addr_hit[48]: begin
        reg_rdata_next[31:0] = hw2reg.data[48].d;
      end

      addr_hit[49]: begin
        reg_rdata_next[31:0] = hw2reg.data[49].d;
      end

      addr_hit[50]: begin
        reg_rdata_next[0] = '0;
      end

      addr_hit[51]: begin
        reg_rdata_next[0] = status_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit))

endmodule

module keccak_reg_top_intf
#(
  parameter int AW = 8,
  localparam int DW = 32
) (
  input logic clk_i,
  input logic rst_ni,
  REG_BUS.in  regbus_slave,
  // To HW
  output keccak_reg_pkg::keccak_reg2hw_t reg2hw, // Write
  input  keccak_reg_pkg::keccak_hw2reg_t hw2reg, // Read
  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);
 localparam int unsigned STRB_WIDTH = DW/8;

`include "register_interface/typedef.svh"
`include "register_interface/assign.svh"

  // Define structs for reg_bus
  typedef logic [AW-1:0] addr_t;
  typedef logic [DW-1:0] data_t;
  typedef logic [STRB_WIDTH-1:0] strb_t;
  `REG_BUS_TYPEDEF_ALL(reg_bus, addr_t, data_t, strb_t)

  reg_bus_req_t s_reg_req;
  reg_bus_rsp_t s_reg_rsp;
  
  // Assign SV interface to structs
  `REG_BUS_ASSIGN_TO_REQ(s_reg_req, regbus_slave)
  `REG_BUS_ASSIGN_FROM_RSP(regbus_slave, s_reg_rsp)

  

  keccak_reg_top #(
    .reg_req_t(reg_bus_req_t),
    .reg_rsp_t(reg_bus_rsp_t),
    .AW(AW)
  ) i_regs (
    .clk_i,
    .rst_ni,
    .reg_req_i(s_reg_req),
    .reg_rsp_o(s_reg_rsp),
    .reg2hw, // Write
    .hw2reg, // Read
    .devmode_i
  );
  
endmodule


