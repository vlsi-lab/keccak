//////////////////////////////////////////////////////////////////////////////////////////
// Authors:      Alessandra Dolmeta - alessandra.dolmeta@polito.it                      //
//               Valeria Piscopo    - valeria.piscopo@polito.it                         //
//               Mattia Mirigaldi    - mattia.mirigaldi@polito.it                       //
// Language:     SystemVerilog                                                          //
// Based on the designed of Michal Peeters and Gilles Van Assche.                       //
//                                                                                      //
//////////////////////////////////////////////////////////////////////////////////////////

// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Top module auto-generated by `reggen`


`include "common_cells/assertions.svh"

module keccak_data_reg_top #(
  parameter type reg_req_t = logic,
  parameter type reg_rsp_t = logic,
  parameter int AW = 9
) (
  input logic clk_i,
  input logic rst_ni,
  input  reg_req_t reg_req_i,
  output reg_rsp_t reg_rsp_o,
  // To HW
  output keccak_data_reg_pkg::keccak_data_reg2hw_t reg2hw, // Write
  input  keccak_data_reg_pkg::keccak_data_hw2reg_t hw2reg, // Read


  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);

  import keccak_data_reg_pkg::* ;

  localparam int DW = 32;
  localparam int DBW = DW/8;                    // Byte Width

  // register signals
  logic           reg_we;
  logic           reg_re;
  logic [AW-1:0]  reg_addr;
  logic [DW-1:0]  reg_wdata;
  logic [DBW-1:0] reg_be;
  logic [DW-1:0]  reg_rdata;
  logic           reg_error;

  logic          addrmiss, wr_err;

  logic [DW-1:0] reg_rdata_next;

  // Below register interface can be changed
  reg_req_t  reg_intf_req;
  reg_rsp_t  reg_intf_rsp;


  assign reg_intf_req = reg_req_i;
  assign reg_rsp_o = reg_intf_rsp;


  assign reg_we = reg_intf_req.valid & reg_intf_req.write;
  assign reg_re = reg_intf_req.valid & ~reg_intf_req.write;
  assign reg_addr = reg_intf_req.addr;
  assign reg_wdata = reg_intf_req.wdata;
  assign reg_be = reg_intf_req.wstrb;
  assign reg_intf_rsp.rdata = reg_rdata;
  assign reg_intf_rsp.error = reg_error;
  assign reg_intf_rsp.ready = 1'b1;

  assign reg_rdata = reg_rdata_next ;
  assign reg_error = (devmode_i & addrmiss) | wr_err;


  // Define SW related signals
  // Format: <reg>_<field>_{wd|we|qs}
  //        or <reg>_{wd|we|qs} if field == 1 or 0
  logic [31:0] din_0_wd;
  logic din_0_we;
  logic [31:0] din_1_wd;
  logic din_1_we;
  logic [31:0] din_2_wd;
  logic din_2_we;
  logic [31:0] din_3_wd;
  logic din_3_we;
  logic [31:0] din_4_wd;
  logic din_4_we;
  logic [31:0] din_5_wd;
  logic din_5_we;
  logic [31:0] din_6_wd;
  logic din_6_we;
  logic [31:0] din_7_wd;
  logic din_7_we;
  logic [31:0] din_8_wd;
  logic din_8_we;
  logic [31:0] din_9_wd;
  logic din_9_we;
  logic [31:0] din_10_wd;
  logic din_10_we;
  logic [31:0] din_11_wd;
  logic din_11_we;
  logic [31:0] din_12_wd;
  logic din_12_we;
  logic [31:0] din_13_wd;
  logic din_13_we;
  logic [31:0] din_14_wd;
  logic din_14_we;
  logic [31:0] din_15_wd;
  logic din_15_we;
  logic [31:0] din_16_wd;
  logic din_16_we;
  logic [31:0] din_17_wd;
  logic din_17_we;
  logic [31:0] din_18_wd;
  logic din_18_we;
  logic [31:0] din_19_wd;
  logic din_19_we;
  logic [31:0] din_20_wd;
  logic din_20_we;
  logic [31:0] din_21_wd;
  logic din_21_we;
  logic [31:0] din_22_wd;
  logic din_22_we;
  logic [31:0] din_23_wd;
  logic din_23_we;
  logic [31:0] din_24_wd;
  logic din_24_we;
  logic [31:0] din_25_wd;
  logic din_25_we;
  logic [31:0] din_26_wd;
  logic din_26_we;
  logic [31:0] din_27_wd;
  logic din_27_we;
  logic [31:0] din_28_wd;
  logic din_28_we;
  logic [31:0] din_29_wd;
  logic din_29_we;
  logic [31:0] din_30_wd;
  logic din_30_we;
  logic [31:0] din_31_wd;
  logic din_31_we;
  logic [31:0] din_32_wd;
  logic din_32_we;
  logic [31:0] din_33_wd;
  logic din_33_we;
  logic [31:0] din_34_wd;
  logic din_34_we;
  logic [31:0] din_35_wd;
  logic din_35_we;
  logic [31:0] din_36_wd;
  logic din_36_we;
  logic [31:0] din_37_wd;
  logic din_37_we;
  logic [31:0] din_38_wd;
  logic din_38_we;
  logic [31:0] din_39_wd;
  logic din_39_we;
  logic [31:0] din_40_wd;
  logic din_40_we;
  logic [31:0] din_41_wd;
  logic din_41_we;
  logic [31:0] din_42_wd;
  logic din_42_we;
  logic [31:0] din_43_wd;
  logic din_43_we;
  logic [31:0] din_44_wd;
  logic din_44_we;
  logic [31:0] din_45_wd;
  logic din_45_we;
  logic [31:0] din_46_wd;
  logic din_46_we;
  logic [31:0] din_47_wd;
  logic din_47_we;
  logic [31:0] din_48_wd;
  logic din_48_we;
  logic [31:0] din_49_wd;
  logic din_49_we;
  logic [31:0] dout_0_qs;
  logic dout_0_re;
  logic [31:0] dout_1_qs;
  logic dout_1_re;
  logic [31:0] dout_2_qs;
  logic dout_2_re;
  logic [31:0] dout_3_qs;
  logic dout_3_re;
  logic [31:0] dout_4_qs;
  logic dout_4_re;
  logic [31:0] dout_5_qs;
  logic dout_5_re;
  logic [31:0] dout_6_qs;
  logic dout_6_re;
  logic [31:0] dout_7_qs;
  logic dout_7_re;
  logic [31:0] dout_8_qs;
  logic dout_8_re;
  logic [31:0] dout_9_qs;
  logic dout_9_re;
  logic [31:0] dout_10_qs;
  logic dout_10_re;
  logic [31:0] dout_11_qs;
  logic dout_11_re;
  logic [31:0] dout_12_qs;
  logic dout_12_re;
  logic [31:0] dout_13_qs;
  logic dout_13_re;
  logic [31:0] dout_14_qs;
  logic dout_14_re;
  logic [31:0] dout_15_qs;
  logic dout_15_re;
  logic [31:0] dout_16_qs;
  logic dout_16_re;
  logic [31:0] dout_17_qs;
  logic dout_17_re;
  logic [31:0] dout_18_qs;
  logic dout_18_re;
  logic [31:0] dout_19_qs;
  logic dout_19_re;
  logic [31:0] dout_20_qs;
  logic dout_20_re;
  logic [31:0] dout_21_qs;
  logic dout_21_re;
  logic [31:0] dout_22_qs;
  logic dout_22_re;
  logic [31:0] dout_23_qs;
  logic dout_23_re;
  logic [31:0] dout_24_qs;
  logic dout_24_re;
  logic [31:0] dout_25_qs;
  logic dout_25_re;
  logic [31:0] dout_26_qs;
  logic dout_26_re;
  logic [31:0] dout_27_qs;
  logic dout_27_re;
  logic [31:0] dout_28_qs;
  logic dout_28_re;
  logic [31:0] dout_29_qs;
  logic dout_29_re;
  logic [31:0] dout_30_qs;
  logic dout_30_re;
  logic [31:0] dout_31_qs;
  logic dout_31_re;
  logic [31:0] dout_32_qs;
  logic dout_32_re;
  logic [31:0] dout_33_qs;
  logic dout_33_re;
  logic [31:0] dout_34_qs;
  logic dout_34_re;
  logic [31:0] dout_35_qs;
  logic dout_35_re;
  logic [31:0] dout_36_qs;
  logic dout_36_re;
  logic [31:0] dout_37_qs;
  logic dout_37_re;
  logic [31:0] dout_38_qs;
  logic dout_38_re;
  logic [31:0] dout_39_qs;
  logic dout_39_re;
  logic [31:0] dout_40_qs;
  logic dout_40_re;
  logic [31:0] dout_41_qs;
  logic dout_41_re;
  logic [31:0] dout_42_qs;
  logic dout_42_re;
  logic [31:0] dout_43_qs;
  logic dout_43_re;
  logic [31:0] dout_44_qs;
  logic dout_44_re;
  logic [31:0] dout_45_qs;
  logic dout_45_re;
  logic [31:0] dout_46_qs;
  logic dout_46_re;
  logic [31:0] dout_47_qs;
  logic dout_47_re;
  logic [31:0] dout_48_qs;
  logic dout_48_re;
  logic [31:0] dout_49_qs;
  logic dout_49_re;

  // Register instances

  // Subregister 0 of Multireg din
  // R[din_0]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_0 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_0_we),
    .wd     (din_0_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[0].q ),

    .qs     ()
  );

  // Subregister 1 of Multireg din
  // R[din_1]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_1 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_1_we),
    .wd     (din_1_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[1].q ),

    .qs     ()
  );

  // Subregister 2 of Multireg din
  // R[din_2]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_2 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_2_we),
    .wd     (din_2_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[2].q ),

    .qs     ()
  );

  // Subregister 3 of Multireg din
  // R[din_3]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_3 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_3_we),
    .wd     (din_3_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[3].q ),

    .qs     ()
  );

  // Subregister 4 of Multireg din
  // R[din_4]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_4 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_4_we),
    .wd     (din_4_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[4].q ),

    .qs     ()
  );

  // Subregister 5 of Multireg din
  // R[din_5]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_5 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_5_we),
    .wd     (din_5_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[5].q ),

    .qs     ()
  );

  // Subregister 6 of Multireg din
  // R[din_6]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_6 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_6_we),
    .wd     (din_6_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[6].q ),

    .qs     ()
  );

  // Subregister 7 of Multireg din
  // R[din_7]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_7 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_7_we),
    .wd     (din_7_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[7].q ),

    .qs     ()
  );

  // Subregister 8 of Multireg din
  // R[din_8]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_8 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_8_we),
    .wd     (din_8_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[8].q ),

    .qs     ()
  );

  // Subregister 9 of Multireg din
  // R[din_9]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_9 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_9_we),
    .wd     (din_9_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[9].q ),

    .qs     ()
  );

  // Subregister 10 of Multireg din
  // R[din_10]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_10 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_10_we),
    .wd     (din_10_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[10].q ),

    .qs     ()
  );

  // Subregister 11 of Multireg din
  // R[din_11]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_11 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_11_we),
    .wd     (din_11_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[11].q ),

    .qs     ()
  );

  // Subregister 12 of Multireg din
  // R[din_12]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_12 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_12_we),
    .wd     (din_12_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[12].q ),

    .qs     ()
  );

  // Subregister 13 of Multireg din
  // R[din_13]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_13 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_13_we),
    .wd     (din_13_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[13].q ),

    .qs     ()
  );

  // Subregister 14 of Multireg din
  // R[din_14]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_14 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_14_we),
    .wd     (din_14_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[14].q ),

    .qs     ()
  );

  // Subregister 15 of Multireg din
  // R[din_15]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_15 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_15_we),
    .wd     (din_15_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[15].q ),

    .qs     ()
  );

  // Subregister 16 of Multireg din
  // R[din_16]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_16 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_16_we),
    .wd     (din_16_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[16].q ),

    .qs     ()
  );

  // Subregister 17 of Multireg din
  // R[din_17]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_17 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_17_we),
    .wd     (din_17_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[17].q ),

    .qs     ()
  );

  // Subregister 18 of Multireg din
  // R[din_18]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_18 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_18_we),
    .wd     (din_18_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[18].q ),

    .qs     ()
  );

  // Subregister 19 of Multireg din
  // R[din_19]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_19 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_19_we),
    .wd     (din_19_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[19].q ),

    .qs     ()
  );

  // Subregister 20 of Multireg din
  // R[din_20]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_20 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_20_we),
    .wd     (din_20_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[20].q ),

    .qs     ()
  );

  // Subregister 21 of Multireg din
  // R[din_21]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_21 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_21_we),
    .wd     (din_21_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[21].q ),

    .qs     ()
  );

  // Subregister 22 of Multireg din
  // R[din_22]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_22 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_22_we),
    .wd     (din_22_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[22].q ),

    .qs     ()
  );

  // Subregister 23 of Multireg din
  // R[din_23]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_23 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_23_we),
    .wd     (din_23_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[23].q ),

    .qs     ()
  );

  // Subregister 24 of Multireg din
  // R[din_24]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_24 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_24_we),
    .wd     (din_24_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[24].q ),

    .qs     ()
  );

  // Subregister 25 of Multireg din
  // R[din_25]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_25 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_25_we),
    .wd     (din_25_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[25].q ),

    .qs     ()
  );

  // Subregister 26 of Multireg din
  // R[din_26]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_26 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_26_we),
    .wd     (din_26_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[26].q ),

    .qs     ()
  );

  // Subregister 27 of Multireg din
  // R[din_27]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_27 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_27_we),
    .wd     (din_27_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[27].q ),

    .qs     ()
  );

  // Subregister 28 of Multireg din
  // R[din_28]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_28 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_28_we),
    .wd     (din_28_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[28].q ),

    .qs     ()
  );

  // Subregister 29 of Multireg din
  // R[din_29]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_29 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_29_we),
    .wd     (din_29_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[29].q ),

    .qs     ()
  );

  // Subregister 30 of Multireg din
  // R[din_30]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_30 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_30_we),
    .wd     (din_30_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[30].q ),

    .qs     ()
  );

  // Subregister 31 of Multireg din
  // R[din_31]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_31 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_31_we),
    .wd     (din_31_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[31].q ),

    .qs     ()
  );

  // Subregister 32 of Multireg din
  // R[din_32]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_32 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_32_we),
    .wd     (din_32_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[32].q ),

    .qs     ()
  );

  // Subregister 33 of Multireg din
  // R[din_33]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_33 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_33_we),
    .wd     (din_33_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[33].q ),

    .qs     ()
  );

  // Subregister 34 of Multireg din
  // R[din_34]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_34 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_34_we),
    .wd     (din_34_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[34].q ),

    .qs     ()
  );

  // Subregister 35 of Multireg din
  // R[din_35]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_35 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_35_we),
    .wd     (din_35_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[35].q ),

    .qs     ()
  );

  // Subregister 36 of Multireg din
  // R[din_36]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_36 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_36_we),
    .wd     (din_36_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[36].q ),

    .qs     ()
  );

  // Subregister 37 of Multireg din
  // R[din_37]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_37 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_37_we),
    .wd     (din_37_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[37].q ),

    .qs     ()
  );

  // Subregister 38 of Multireg din
  // R[din_38]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_38 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_38_we),
    .wd     (din_38_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[38].q ),

    .qs     ()
  );

  // Subregister 39 of Multireg din
  // R[din_39]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_39 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_39_we),
    .wd     (din_39_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[39].q ),

    .qs     ()
  );

  // Subregister 40 of Multireg din
  // R[din_40]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_40 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_40_we),
    .wd     (din_40_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[40].q ),

    .qs     ()
  );

  // Subregister 41 of Multireg din
  // R[din_41]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_41 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_41_we),
    .wd     (din_41_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[41].q ),

    .qs     ()
  );

  // Subregister 42 of Multireg din
  // R[din_42]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_42 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_42_we),
    .wd     (din_42_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[42].q ),

    .qs     ()
  );

  // Subregister 43 of Multireg din
  // R[din_43]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_43 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_43_we),
    .wd     (din_43_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[43].q ),

    .qs     ()
  );

  // Subregister 44 of Multireg din
  // R[din_44]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_44 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_44_we),
    .wd     (din_44_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[44].q ),

    .qs     ()
  );

  // Subregister 45 of Multireg din
  // R[din_45]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_45 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_45_we),
    .wd     (din_45_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[45].q ),

    .qs     ()
  );

  // Subregister 46 of Multireg din
  // R[din_46]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_46 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_46_we),
    .wd     (din_46_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[46].q ),

    .qs     ()
  );

  // Subregister 47 of Multireg din
  // R[din_47]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_47 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_47_we),
    .wd     (din_47_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[47].q ),

    .qs     ()
  );

  // Subregister 48 of Multireg din
  // R[din_48]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_48 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_48_we),
    .wd     (din_48_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[48].q ),

    .qs     ()
  );

  // Subregister 49 of Multireg din
  // R[din_49]: V(False)

  prim_subreg #(
    .DW      (32),
    .SWACCESS("WO"),
    .RESVAL  (32'h0)
  ) u_din_49 (
    .clk_i   (clk_i    ),
    .rst_ni  (rst_ni  ),

    // from register interface
    .we     (din_49_we),
    .wd     (din_49_wd),

    // from internal hardware
    .de     (1'b0),
    .d      ('0  ),

    // to internal hardware
    .qe     (),
    .q      (reg2hw.din[49].q ),

    .qs     ()
  );



  // Subregister 0 of Multireg dout
  // R[dout_0]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_0 (
    .re     (dout_0_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[0].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_0_qs)
  );

  // Subregister 1 of Multireg dout
  // R[dout_1]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_1 (
    .re     (dout_1_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[1].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_1_qs)
  );

  // Subregister 2 of Multireg dout
  // R[dout_2]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_2 (
    .re     (dout_2_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[2].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_2_qs)
  );

  // Subregister 3 of Multireg dout
  // R[dout_3]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_3 (
    .re     (dout_3_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[3].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_3_qs)
  );

  // Subregister 4 of Multireg dout
  // R[dout_4]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_4 (
    .re     (dout_4_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[4].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_4_qs)
  );

  // Subregister 5 of Multireg dout
  // R[dout_5]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_5 (
    .re     (dout_5_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[5].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_5_qs)
  );

  // Subregister 6 of Multireg dout
  // R[dout_6]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_6 (
    .re     (dout_6_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[6].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_6_qs)
  );

  // Subregister 7 of Multireg dout
  // R[dout_7]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_7 (
    .re     (dout_7_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[7].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_7_qs)
  );

  // Subregister 8 of Multireg dout
  // R[dout_8]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_8 (
    .re     (dout_8_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[8].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_8_qs)
  );

  // Subregister 9 of Multireg dout
  // R[dout_9]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_9 (
    .re     (dout_9_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[9].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_9_qs)
  );

  // Subregister 10 of Multireg dout
  // R[dout_10]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_10 (
    .re     (dout_10_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[10].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_10_qs)
  );

  // Subregister 11 of Multireg dout
  // R[dout_11]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_11 (
    .re     (dout_11_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[11].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_11_qs)
  );

  // Subregister 12 of Multireg dout
  // R[dout_12]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_12 (
    .re     (dout_12_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[12].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_12_qs)
  );

  // Subregister 13 of Multireg dout
  // R[dout_13]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_13 (
    .re     (dout_13_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[13].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_13_qs)
  );

  // Subregister 14 of Multireg dout
  // R[dout_14]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_14 (
    .re     (dout_14_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[14].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_14_qs)
  );

  // Subregister 15 of Multireg dout
  // R[dout_15]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_15 (
    .re     (dout_15_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[15].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_15_qs)
  );

  // Subregister 16 of Multireg dout
  // R[dout_16]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_16 (
    .re     (dout_16_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[16].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_16_qs)
  );

  // Subregister 17 of Multireg dout
  // R[dout_17]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_17 (
    .re     (dout_17_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[17].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_17_qs)
  );

  // Subregister 18 of Multireg dout
  // R[dout_18]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_18 (
    .re     (dout_18_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[18].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_18_qs)
  );

  // Subregister 19 of Multireg dout
  // R[dout_19]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_19 (
    .re     (dout_19_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[19].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_19_qs)
  );

  // Subregister 20 of Multireg dout
  // R[dout_20]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_20 (
    .re     (dout_20_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[20].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_20_qs)
  );

  // Subregister 21 of Multireg dout
  // R[dout_21]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_21 (
    .re     (dout_21_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[21].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_21_qs)
  );

  // Subregister 22 of Multireg dout
  // R[dout_22]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_22 (
    .re     (dout_22_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[22].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_22_qs)
  );

  // Subregister 23 of Multireg dout
  // R[dout_23]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_23 (
    .re     (dout_23_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[23].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_23_qs)
  );

  // Subregister 24 of Multireg dout
  // R[dout_24]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_24 (
    .re     (dout_24_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[24].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_24_qs)
  );

  // Subregister 25 of Multireg dout
  // R[dout_25]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_25 (
    .re     (dout_25_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[25].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_25_qs)
  );

  // Subregister 26 of Multireg dout
  // R[dout_26]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_26 (
    .re     (dout_26_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[26].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_26_qs)
  );

  // Subregister 27 of Multireg dout
  // R[dout_27]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_27 (
    .re     (dout_27_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[27].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_27_qs)
  );

  // Subregister 28 of Multireg dout
  // R[dout_28]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_28 (
    .re     (dout_28_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[28].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_28_qs)
  );

  // Subregister 29 of Multireg dout
  // R[dout_29]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_29 (
    .re     (dout_29_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[29].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_29_qs)
  );

  // Subregister 30 of Multireg dout
  // R[dout_30]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_30 (
    .re     (dout_30_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[30].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_30_qs)
  );

  // Subregister 31 of Multireg dout
  // R[dout_31]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_31 (
    .re     (dout_31_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[31].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_31_qs)
  );

  // Subregister 32 of Multireg dout
  // R[dout_32]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_32 (
    .re     (dout_32_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[32].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_32_qs)
  );

  // Subregister 33 of Multireg dout
  // R[dout_33]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_33 (
    .re     (dout_33_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[33].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_33_qs)
  );

  // Subregister 34 of Multireg dout
  // R[dout_34]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_34 (
    .re     (dout_34_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[34].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_34_qs)
  );

  // Subregister 35 of Multireg dout
  // R[dout_35]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_35 (
    .re     (dout_35_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[35].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_35_qs)
  );

  // Subregister 36 of Multireg dout
  // R[dout_36]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_36 (
    .re     (dout_36_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[36].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_36_qs)
  );

  // Subregister 37 of Multireg dout
  // R[dout_37]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_37 (
    .re     (dout_37_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[37].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_37_qs)
  );

  // Subregister 38 of Multireg dout
  // R[dout_38]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_38 (
    .re     (dout_38_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[38].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_38_qs)
  );

  // Subregister 39 of Multireg dout
  // R[dout_39]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_39 (
    .re     (dout_39_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[39].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_39_qs)
  );

  // Subregister 40 of Multireg dout
  // R[dout_40]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_40 (
    .re     (dout_40_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[40].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_40_qs)
  );

  // Subregister 41 of Multireg dout
  // R[dout_41]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_41 (
    .re     (dout_41_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[41].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_41_qs)
  );

  // Subregister 42 of Multireg dout
  // R[dout_42]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_42 (
    .re     (dout_42_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[42].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_42_qs)
  );

  // Subregister 43 of Multireg dout
  // R[dout_43]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_43 (
    .re     (dout_43_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[43].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_43_qs)
  );

  // Subregister 44 of Multireg dout
  // R[dout_44]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_44 (
    .re     (dout_44_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[44].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_44_qs)
  );

  // Subregister 45 of Multireg dout
  // R[dout_45]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_45 (
    .re     (dout_45_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[45].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_45_qs)
  );

  // Subregister 46 of Multireg dout
  // R[dout_46]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_46 (
    .re     (dout_46_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[46].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_46_qs)
  );

  // Subregister 47 of Multireg dout
  // R[dout_47]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_47 (
    .re     (dout_47_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[47].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_47_qs)
  );

  // Subregister 48 of Multireg dout
  // R[dout_48]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_48 (
    .re     (dout_48_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[48].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_48_qs)
  );

  // Subregister 49 of Multireg dout
  // R[dout_49]: V(True)

  prim_subreg_ext #(
    .DW    (32)
  ) u_dout_49 (
    .re     (dout_49_re),
    .we     (1'b0),
    .wd     ('0),
    .d      (hw2reg.dout[49].d),
    .qre    (),
    .qe     (),
    .q      (),
    .qs     (dout_49_qs)
  );




  logic [99:0] addr_hit;
  always_comb begin
    addr_hit = '0;
    addr_hit[ 0] = (reg_addr == KECCAK_DATA_DIN_0_OFFSET);
    addr_hit[ 1] = (reg_addr == KECCAK_DATA_DIN_1_OFFSET);
    addr_hit[ 2] = (reg_addr == KECCAK_DATA_DIN_2_OFFSET);
    addr_hit[ 3] = (reg_addr == KECCAK_DATA_DIN_3_OFFSET);
    addr_hit[ 4] = (reg_addr == KECCAK_DATA_DIN_4_OFFSET);
    addr_hit[ 5] = (reg_addr == KECCAK_DATA_DIN_5_OFFSET);
    addr_hit[ 6] = (reg_addr == KECCAK_DATA_DIN_6_OFFSET);
    addr_hit[ 7] = (reg_addr == KECCAK_DATA_DIN_7_OFFSET);
    addr_hit[ 8] = (reg_addr == KECCAK_DATA_DIN_8_OFFSET);
    addr_hit[ 9] = (reg_addr == KECCAK_DATA_DIN_9_OFFSET);
    addr_hit[10] = (reg_addr == KECCAK_DATA_DIN_10_OFFSET);
    addr_hit[11] = (reg_addr == KECCAK_DATA_DIN_11_OFFSET);
    addr_hit[12] = (reg_addr == KECCAK_DATA_DIN_12_OFFSET);
    addr_hit[13] = (reg_addr == KECCAK_DATA_DIN_13_OFFSET);
    addr_hit[14] = (reg_addr == KECCAK_DATA_DIN_14_OFFSET);
    addr_hit[15] = (reg_addr == KECCAK_DATA_DIN_15_OFFSET);
    addr_hit[16] = (reg_addr == KECCAK_DATA_DIN_16_OFFSET);
    addr_hit[17] = (reg_addr == KECCAK_DATA_DIN_17_OFFSET);
    addr_hit[18] = (reg_addr == KECCAK_DATA_DIN_18_OFFSET);
    addr_hit[19] = (reg_addr == KECCAK_DATA_DIN_19_OFFSET);
    addr_hit[20] = (reg_addr == KECCAK_DATA_DIN_20_OFFSET);
    addr_hit[21] = (reg_addr == KECCAK_DATA_DIN_21_OFFSET);
    addr_hit[22] = (reg_addr == KECCAK_DATA_DIN_22_OFFSET);
    addr_hit[23] = (reg_addr == KECCAK_DATA_DIN_23_OFFSET);
    addr_hit[24] = (reg_addr == KECCAK_DATA_DIN_24_OFFSET);
    addr_hit[25] = (reg_addr == KECCAK_DATA_DIN_25_OFFSET);
    addr_hit[26] = (reg_addr == KECCAK_DATA_DIN_26_OFFSET);
    addr_hit[27] = (reg_addr == KECCAK_DATA_DIN_27_OFFSET);
    addr_hit[28] = (reg_addr == KECCAK_DATA_DIN_28_OFFSET);
    addr_hit[29] = (reg_addr == KECCAK_DATA_DIN_29_OFFSET);
    addr_hit[30] = (reg_addr == KECCAK_DATA_DIN_30_OFFSET);
    addr_hit[31] = (reg_addr == KECCAK_DATA_DIN_31_OFFSET);
    addr_hit[32] = (reg_addr == KECCAK_DATA_DIN_32_OFFSET);
    addr_hit[33] = (reg_addr == KECCAK_DATA_DIN_33_OFFSET);
    addr_hit[34] = (reg_addr == KECCAK_DATA_DIN_34_OFFSET);
    addr_hit[35] = (reg_addr == KECCAK_DATA_DIN_35_OFFSET);
    addr_hit[36] = (reg_addr == KECCAK_DATA_DIN_36_OFFSET);
    addr_hit[37] = (reg_addr == KECCAK_DATA_DIN_37_OFFSET);
    addr_hit[38] = (reg_addr == KECCAK_DATA_DIN_38_OFFSET);
    addr_hit[39] = (reg_addr == KECCAK_DATA_DIN_39_OFFSET);
    addr_hit[40] = (reg_addr == KECCAK_DATA_DIN_40_OFFSET);
    addr_hit[41] = (reg_addr == KECCAK_DATA_DIN_41_OFFSET);
    addr_hit[42] = (reg_addr == KECCAK_DATA_DIN_42_OFFSET);
    addr_hit[43] = (reg_addr == KECCAK_DATA_DIN_43_OFFSET);
    addr_hit[44] = (reg_addr == KECCAK_DATA_DIN_44_OFFSET);
    addr_hit[45] = (reg_addr == KECCAK_DATA_DIN_45_OFFSET);
    addr_hit[46] = (reg_addr == KECCAK_DATA_DIN_46_OFFSET);
    addr_hit[47] = (reg_addr == KECCAK_DATA_DIN_47_OFFSET);
    addr_hit[48] = (reg_addr == KECCAK_DATA_DIN_48_OFFSET);
    addr_hit[49] = (reg_addr == KECCAK_DATA_DIN_49_OFFSET);
    addr_hit[50] = (reg_addr == KECCAK_DATA_DOUT_0_OFFSET);
    addr_hit[51] = (reg_addr == KECCAK_DATA_DOUT_1_OFFSET);
    addr_hit[52] = (reg_addr == KECCAK_DATA_DOUT_2_OFFSET);
    addr_hit[53] = (reg_addr == KECCAK_DATA_DOUT_3_OFFSET);
    addr_hit[54] = (reg_addr == KECCAK_DATA_DOUT_4_OFFSET);
    addr_hit[55] = (reg_addr == KECCAK_DATA_DOUT_5_OFFSET);
    addr_hit[56] = (reg_addr == KECCAK_DATA_DOUT_6_OFFSET);
    addr_hit[57] = (reg_addr == KECCAK_DATA_DOUT_7_OFFSET);
    addr_hit[58] = (reg_addr == KECCAK_DATA_DOUT_8_OFFSET);
    addr_hit[59] = (reg_addr == KECCAK_DATA_DOUT_9_OFFSET);
    addr_hit[60] = (reg_addr == KECCAK_DATA_DOUT_10_OFFSET);
    addr_hit[61] = (reg_addr == KECCAK_DATA_DOUT_11_OFFSET);
    addr_hit[62] = (reg_addr == KECCAK_DATA_DOUT_12_OFFSET);
    addr_hit[63] = (reg_addr == KECCAK_DATA_DOUT_13_OFFSET);
    addr_hit[64] = (reg_addr == KECCAK_DATA_DOUT_14_OFFSET);
    addr_hit[65] = (reg_addr == KECCAK_DATA_DOUT_15_OFFSET);
    addr_hit[66] = (reg_addr == KECCAK_DATA_DOUT_16_OFFSET);
    addr_hit[67] = (reg_addr == KECCAK_DATA_DOUT_17_OFFSET);
    addr_hit[68] = (reg_addr == KECCAK_DATA_DOUT_18_OFFSET);
    addr_hit[69] = (reg_addr == KECCAK_DATA_DOUT_19_OFFSET);
    addr_hit[70] = (reg_addr == KECCAK_DATA_DOUT_20_OFFSET);
    addr_hit[71] = (reg_addr == KECCAK_DATA_DOUT_21_OFFSET);
    addr_hit[72] = (reg_addr == KECCAK_DATA_DOUT_22_OFFSET);
    addr_hit[73] = (reg_addr == KECCAK_DATA_DOUT_23_OFFSET);
    addr_hit[74] = (reg_addr == KECCAK_DATA_DOUT_24_OFFSET);
    addr_hit[75] = (reg_addr == KECCAK_DATA_DOUT_25_OFFSET);
    addr_hit[76] = (reg_addr == KECCAK_DATA_DOUT_26_OFFSET);
    addr_hit[77] = (reg_addr == KECCAK_DATA_DOUT_27_OFFSET);
    addr_hit[78] = (reg_addr == KECCAK_DATA_DOUT_28_OFFSET);
    addr_hit[79] = (reg_addr == KECCAK_DATA_DOUT_29_OFFSET);
    addr_hit[80] = (reg_addr == KECCAK_DATA_DOUT_30_OFFSET);
    addr_hit[81] = (reg_addr == KECCAK_DATA_DOUT_31_OFFSET);
    addr_hit[82] = (reg_addr == KECCAK_DATA_DOUT_32_OFFSET);
    addr_hit[83] = (reg_addr == KECCAK_DATA_DOUT_33_OFFSET);
    addr_hit[84] = (reg_addr == KECCAK_DATA_DOUT_34_OFFSET);
    addr_hit[85] = (reg_addr == KECCAK_DATA_DOUT_35_OFFSET);
    addr_hit[86] = (reg_addr == KECCAK_DATA_DOUT_36_OFFSET);
    addr_hit[87] = (reg_addr == KECCAK_DATA_DOUT_37_OFFSET);
    addr_hit[88] = (reg_addr == KECCAK_DATA_DOUT_38_OFFSET);
    addr_hit[89] = (reg_addr == KECCAK_DATA_DOUT_39_OFFSET);
    addr_hit[90] = (reg_addr == KECCAK_DATA_DOUT_40_OFFSET);
    addr_hit[91] = (reg_addr == KECCAK_DATA_DOUT_41_OFFSET);
    addr_hit[92] = (reg_addr == KECCAK_DATA_DOUT_42_OFFSET);
    addr_hit[93] = (reg_addr == KECCAK_DATA_DOUT_43_OFFSET);
    addr_hit[94] = (reg_addr == KECCAK_DATA_DOUT_44_OFFSET);
    addr_hit[95] = (reg_addr == KECCAK_DATA_DOUT_45_OFFSET);
    addr_hit[96] = (reg_addr == KECCAK_DATA_DOUT_46_OFFSET);
    addr_hit[97] = (reg_addr == KECCAK_DATA_DOUT_47_OFFSET);
    addr_hit[98] = (reg_addr == KECCAK_DATA_DOUT_48_OFFSET);
    addr_hit[99] = (reg_addr == KECCAK_DATA_DOUT_49_OFFSET);
  end

  assign addrmiss = (reg_re || reg_we) ? ~|addr_hit : 1'b0 ;

  // Check sub-word write is permitted
  always_comb begin
    wr_err = (reg_we &
              ((addr_hit[ 0] & (|(KECCAK_DATA_PERMIT[ 0] & ~reg_be))) |
               (addr_hit[ 1] & (|(KECCAK_DATA_PERMIT[ 1] & ~reg_be))) |
               (addr_hit[ 2] & (|(KECCAK_DATA_PERMIT[ 2] & ~reg_be))) |
               (addr_hit[ 3] & (|(KECCAK_DATA_PERMIT[ 3] & ~reg_be))) |
               (addr_hit[ 4] & (|(KECCAK_DATA_PERMIT[ 4] & ~reg_be))) |
               (addr_hit[ 5] & (|(KECCAK_DATA_PERMIT[ 5] & ~reg_be))) |
               (addr_hit[ 6] & (|(KECCAK_DATA_PERMIT[ 6] & ~reg_be))) |
               (addr_hit[ 7] & (|(KECCAK_DATA_PERMIT[ 7] & ~reg_be))) |
               (addr_hit[ 8] & (|(KECCAK_DATA_PERMIT[ 8] & ~reg_be))) |
               (addr_hit[ 9] & (|(KECCAK_DATA_PERMIT[ 9] & ~reg_be))) |
               (addr_hit[10] & (|(KECCAK_DATA_PERMIT[10] & ~reg_be))) |
               (addr_hit[11] & (|(KECCAK_DATA_PERMIT[11] & ~reg_be))) |
               (addr_hit[12] & (|(KECCAK_DATA_PERMIT[12] & ~reg_be))) |
               (addr_hit[13] & (|(KECCAK_DATA_PERMIT[13] & ~reg_be))) |
               (addr_hit[14] & (|(KECCAK_DATA_PERMIT[14] & ~reg_be))) |
               (addr_hit[15] & (|(KECCAK_DATA_PERMIT[15] & ~reg_be))) |
               (addr_hit[16] & (|(KECCAK_DATA_PERMIT[16] & ~reg_be))) |
               (addr_hit[17] & (|(KECCAK_DATA_PERMIT[17] & ~reg_be))) |
               (addr_hit[18] & (|(KECCAK_DATA_PERMIT[18] & ~reg_be))) |
               (addr_hit[19] & (|(KECCAK_DATA_PERMIT[19] & ~reg_be))) |
               (addr_hit[20] & (|(KECCAK_DATA_PERMIT[20] & ~reg_be))) |
               (addr_hit[21] & (|(KECCAK_DATA_PERMIT[21] & ~reg_be))) |
               (addr_hit[22] & (|(KECCAK_DATA_PERMIT[22] & ~reg_be))) |
               (addr_hit[23] & (|(KECCAK_DATA_PERMIT[23] & ~reg_be))) |
               (addr_hit[24] & (|(KECCAK_DATA_PERMIT[24] & ~reg_be))) |
               (addr_hit[25] & (|(KECCAK_DATA_PERMIT[25] & ~reg_be))) |
               (addr_hit[26] & (|(KECCAK_DATA_PERMIT[26] & ~reg_be))) |
               (addr_hit[27] & (|(KECCAK_DATA_PERMIT[27] & ~reg_be))) |
               (addr_hit[28] & (|(KECCAK_DATA_PERMIT[28] & ~reg_be))) |
               (addr_hit[29] & (|(KECCAK_DATA_PERMIT[29] & ~reg_be))) |
               (addr_hit[30] & (|(KECCAK_DATA_PERMIT[30] & ~reg_be))) |
               (addr_hit[31] & (|(KECCAK_DATA_PERMIT[31] & ~reg_be))) |
               (addr_hit[32] & (|(KECCAK_DATA_PERMIT[32] & ~reg_be))) |
               (addr_hit[33] & (|(KECCAK_DATA_PERMIT[33] & ~reg_be))) |
               (addr_hit[34] & (|(KECCAK_DATA_PERMIT[34] & ~reg_be))) |
               (addr_hit[35] & (|(KECCAK_DATA_PERMIT[35] & ~reg_be))) |
               (addr_hit[36] & (|(KECCAK_DATA_PERMIT[36] & ~reg_be))) |
               (addr_hit[37] & (|(KECCAK_DATA_PERMIT[37] & ~reg_be))) |
               (addr_hit[38] & (|(KECCAK_DATA_PERMIT[38] & ~reg_be))) |
               (addr_hit[39] & (|(KECCAK_DATA_PERMIT[39] & ~reg_be))) |
               (addr_hit[40] & (|(KECCAK_DATA_PERMIT[40] & ~reg_be))) |
               (addr_hit[41] & (|(KECCAK_DATA_PERMIT[41] & ~reg_be))) |
               (addr_hit[42] & (|(KECCAK_DATA_PERMIT[42] & ~reg_be))) |
               (addr_hit[43] & (|(KECCAK_DATA_PERMIT[43] & ~reg_be))) |
               (addr_hit[44] & (|(KECCAK_DATA_PERMIT[44] & ~reg_be))) |
               (addr_hit[45] & (|(KECCAK_DATA_PERMIT[45] & ~reg_be))) |
               (addr_hit[46] & (|(KECCAK_DATA_PERMIT[46] & ~reg_be))) |
               (addr_hit[47] & (|(KECCAK_DATA_PERMIT[47] & ~reg_be))) |
               (addr_hit[48] & (|(KECCAK_DATA_PERMIT[48] & ~reg_be))) |
               (addr_hit[49] & (|(KECCAK_DATA_PERMIT[49] & ~reg_be))) |
               (addr_hit[50] & (|(KECCAK_DATA_PERMIT[50] & ~reg_be))) |
               (addr_hit[51] & (|(KECCAK_DATA_PERMIT[51] & ~reg_be))) |
               (addr_hit[52] & (|(KECCAK_DATA_PERMIT[52] & ~reg_be))) |
               (addr_hit[53] & (|(KECCAK_DATA_PERMIT[53] & ~reg_be))) |
               (addr_hit[54] & (|(KECCAK_DATA_PERMIT[54] & ~reg_be))) |
               (addr_hit[55] & (|(KECCAK_DATA_PERMIT[55] & ~reg_be))) |
               (addr_hit[56] & (|(KECCAK_DATA_PERMIT[56] & ~reg_be))) |
               (addr_hit[57] & (|(KECCAK_DATA_PERMIT[57] & ~reg_be))) |
               (addr_hit[58] & (|(KECCAK_DATA_PERMIT[58] & ~reg_be))) |
               (addr_hit[59] & (|(KECCAK_DATA_PERMIT[59] & ~reg_be))) |
               (addr_hit[60] & (|(KECCAK_DATA_PERMIT[60] & ~reg_be))) |
               (addr_hit[61] & (|(KECCAK_DATA_PERMIT[61] & ~reg_be))) |
               (addr_hit[62] & (|(KECCAK_DATA_PERMIT[62] & ~reg_be))) |
               (addr_hit[63] & (|(KECCAK_DATA_PERMIT[63] & ~reg_be))) |
               (addr_hit[64] & (|(KECCAK_DATA_PERMIT[64] & ~reg_be))) |
               (addr_hit[65] & (|(KECCAK_DATA_PERMIT[65] & ~reg_be))) |
               (addr_hit[66] & (|(KECCAK_DATA_PERMIT[66] & ~reg_be))) |
               (addr_hit[67] & (|(KECCAK_DATA_PERMIT[67] & ~reg_be))) |
               (addr_hit[68] & (|(KECCAK_DATA_PERMIT[68] & ~reg_be))) |
               (addr_hit[69] & (|(KECCAK_DATA_PERMIT[69] & ~reg_be))) |
               (addr_hit[70] & (|(KECCAK_DATA_PERMIT[70] & ~reg_be))) |
               (addr_hit[71] & (|(KECCAK_DATA_PERMIT[71] & ~reg_be))) |
               (addr_hit[72] & (|(KECCAK_DATA_PERMIT[72] & ~reg_be))) |
               (addr_hit[73] & (|(KECCAK_DATA_PERMIT[73] & ~reg_be))) |
               (addr_hit[74] & (|(KECCAK_DATA_PERMIT[74] & ~reg_be))) |
               (addr_hit[75] & (|(KECCAK_DATA_PERMIT[75] & ~reg_be))) |
               (addr_hit[76] & (|(KECCAK_DATA_PERMIT[76] & ~reg_be))) |
               (addr_hit[77] & (|(KECCAK_DATA_PERMIT[77] & ~reg_be))) |
               (addr_hit[78] & (|(KECCAK_DATA_PERMIT[78] & ~reg_be))) |
               (addr_hit[79] & (|(KECCAK_DATA_PERMIT[79] & ~reg_be))) |
               (addr_hit[80] & (|(KECCAK_DATA_PERMIT[80] & ~reg_be))) |
               (addr_hit[81] & (|(KECCAK_DATA_PERMIT[81] & ~reg_be))) |
               (addr_hit[82] & (|(KECCAK_DATA_PERMIT[82] & ~reg_be))) |
               (addr_hit[83] & (|(KECCAK_DATA_PERMIT[83] & ~reg_be))) |
               (addr_hit[84] & (|(KECCAK_DATA_PERMIT[84] & ~reg_be))) |
               (addr_hit[85] & (|(KECCAK_DATA_PERMIT[85] & ~reg_be))) |
               (addr_hit[86] & (|(KECCAK_DATA_PERMIT[86] & ~reg_be))) |
               (addr_hit[87] & (|(KECCAK_DATA_PERMIT[87] & ~reg_be))) |
               (addr_hit[88] & (|(KECCAK_DATA_PERMIT[88] & ~reg_be))) |
               (addr_hit[89] & (|(KECCAK_DATA_PERMIT[89] & ~reg_be))) |
               (addr_hit[90] & (|(KECCAK_DATA_PERMIT[90] & ~reg_be))) |
               (addr_hit[91] & (|(KECCAK_DATA_PERMIT[91] & ~reg_be))) |
               (addr_hit[92] & (|(KECCAK_DATA_PERMIT[92] & ~reg_be))) |
               (addr_hit[93] & (|(KECCAK_DATA_PERMIT[93] & ~reg_be))) |
               (addr_hit[94] & (|(KECCAK_DATA_PERMIT[94] & ~reg_be))) |
               (addr_hit[95] & (|(KECCAK_DATA_PERMIT[95] & ~reg_be))) |
               (addr_hit[96] & (|(KECCAK_DATA_PERMIT[96] & ~reg_be))) |
               (addr_hit[97] & (|(KECCAK_DATA_PERMIT[97] & ~reg_be))) |
               (addr_hit[98] & (|(KECCAK_DATA_PERMIT[98] & ~reg_be))) |
               (addr_hit[99] & (|(KECCAK_DATA_PERMIT[99] & ~reg_be)))));
  end

  assign din_0_we = addr_hit[0] & reg_we & !reg_error;
  assign din_0_wd = reg_wdata[31:0];

  assign din_1_we = addr_hit[1] & reg_we & !reg_error;
  assign din_1_wd = reg_wdata[31:0];

  assign din_2_we = addr_hit[2] & reg_we & !reg_error;
  assign din_2_wd = reg_wdata[31:0];

  assign din_3_we = addr_hit[3] & reg_we & !reg_error;
  assign din_3_wd = reg_wdata[31:0];

  assign din_4_we = addr_hit[4] & reg_we & !reg_error;
  assign din_4_wd = reg_wdata[31:0];

  assign din_5_we = addr_hit[5] & reg_we & !reg_error;
  assign din_5_wd = reg_wdata[31:0];

  assign din_6_we = addr_hit[6] & reg_we & !reg_error;
  assign din_6_wd = reg_wdata[31:0];

  assign din_7_we = addr_hit[7] & reg_we & !reg_error;
  assign din_7_wd = reg_wdata[31:0];

  assign din_8_we = addr_hit[8] & reg_we & !reg_error;
  assign din_8_wd = reg_wdata[31:0];

  assign din_9_we = addr_hit[9] & reg_we & !reg_error;
  assign din_9_wd = reg_wdata[31:0];

  assign din_10_we = addr_hit[10] & reg_we & !reg_error;
  assign din_10_wd = reg_wdata[31:0];

  assign din_11_we = addr_hit[11] & reg_we & !reg_error;
  assign din_11_wd = reg_wdata[31:0];

  assign din_12_we = addr_hit[12] & reg_we & !reg_error;
  assign din_12_wd = reg_wdata[31:0];

  assign din_13_we = addr_hit[13] & reg_we & !reg_error;
  assign din_13_wd = reg_wdata[31:0];

  assign din_14_we = addr_hit[14] & reg_we & !reg_error;
  assign din_14_wd = reg_wdata[31:0];

  assign din_15_we = addr_hit[15] & reg_we & !reg_error;
  assign din_15_wd = reg_wdata[31:0];

  assign din_16_we = addr_hit[16] & reg_we & !reg_error;
  assign din_16_wd = reg_wdata[31:0];

  assign din_17_we = addr_hit[17] & reg_we & !reg_error;
  assign din_17_wd = reg_wdata[31:0];

  assign din_18_we = addr_hit[18] & reg_we & !reg_error;
  assign din_18_wd = reg_wdata[31:0];

  assign din_19_we = addr_hit[19] & reg_we & !reg_error;
  assign din_19_wd = reg_wdata[31:0];

  assign din_20_we = addr_hit[20] & reg_we & !reg_error;
  assign din_20_wd = reg_wdata[31:0];

  assign din_21_we = addr_hit[21] & reg_we & !reg_error;
  assign din_21_wd = reg_wdata[31:0];

  assign din_22_we = addr_hit[22] & reg_we & !reg_error;
  assign din_22_wd = reg_wdata[31:0];

  assign din_23_we = addr_hit[23] & reg_we & !reg_error;
  assign din_23_wd = reg_wdata[31:0];

  assign din_24_we = addr_hit[24] & reg_we & !reg_error;
  assign din_24_wd = reg_wdata[31:0];

  assign din_25_we = addr_hit[25] & reg_we & !reg_error;
  assign din_25_wd = reg_wdata[31:0];

  assign din_26_we = addr_hit[26] & reg_we & !reg_error;
  assign din_26_wd = reg_wdata[31:0];

  assign din_27_we = addr_hit[27] & reg_we & !reg_error;
  assign din_27_wd = reg_wdata[31:0];

  assign din_28_we = addr_hit[28] & reg_we & !reg_error;
  assign din_28_wd = reg_wdata[31:0];

  assign din_29_we = addr_hit[29] & reg_we & !reg_error;
  assign din_29_wd = reg_wdata[31:0];

  assign din_30_we = addr_hit[30] & reg_we & !reg_error;
  assign din_30_wd = reg_wdata[31:0];

  assign din_31_we = addr_hit[31] & reg_we & !reg_error;
  assign din_31_wd = reg_wdata[31:0];

  assign din_32_we = addr_hit[32] & reg_we & !reg_error;
  assign din_32_wd = reg_wdata[31:0];

  assign din_33_we = addr_hit[33] & reg_we & !reg_error;
  assign din_33_wd = reg_wdata[31:0];

  assign din_34_we = addr_hit[34] & reg_we & !reg_error;
  assign din_34_wd = reg_wdata[31:0];

  assign din_35_we = addr_hit[35] & reg_we & !reg_error;
  assign din_35_wd = reg_wdata[31:0];

  assign din_36_we = addr_hit[36] & reg_we & !reg_error;
  assign din_36_wd = reg_wdata[31:0];

  assign din_37_we = addr_hit[37] & reg_we & !reg_error;
  assign din_37_wd = reg_wdata[31:0];

  assign din_38_we = addr_hit[38] & reg_we & !reg_error;
  assign din_38_wd = reg_wdata[31:0];

  assign din_39_we = addr_hit[39] & reg_we & !reg_error;
  assign din_39_wd = reg_wdata[31:0];

  assign din_40_we = addr_hit[40] & reg_we & !reg_error;
  assign din_40_wd = reg_wdata[31:0];

  assign din_41_we = addr_hit[41] & reg_we & !reg_error;
  assign din_41_wd = reg_wdata[31:0];

  assign din_42_we = addr_hit[42] & reg_we & !reg_error;
  assign din_42_wd = reg_wdata[31:0];

  assign din_43_we = addr_hit[43] & reg_we & !reg_error;
  assign din_43_wd = reg_wdata[31:0];

  assign din_44_we = addr_hit[44] & reg_we & !reg_error;
  assign din_44_wd = reg_wdata[31:0];

  assign din_45_we = addr_hit[45] & reg_we & !reg_error;
  assign din_45_wd = reg_wdata[31:0];

  assign din_46_we = addr_hit[46] & reg_we & !reg_error;
  assign din_46_wd = reg_wdata[31:0];

  assign din_47_we = addr_hit[47] & reg_we & !reg_error;
  assign din_47_wd = reg_wdata[31:0];

  assign din_48_we = addr_hit[48] & reg_we & !reg_error;
  assign din_48_wd = reg_wdata[31:0];

  assign din_49_we = addr_hit[49] & reg_we & !reg_error;
  assign din_49_wd = reg_wdata[31:0];

  assign dout_0_re = addr_hit[50] & reg_re & !reg_error;

  assign dout_1_re = addr_hit[51] & reg_re & !reg_error;

  assign dout_2_re = addr_hit[52] & reg_re & !reg_error;

  assign dout_3_re = addr_hit[53] & reg_re & !reg_error;

  assign dout_4_re = addr_hit[54] & reg_re & !reg_error;

  assign dout_5_re = addr_hit[55] & reg_re & !reg_error;

  assign dout_6_re = addr_hit[56] & reg_re & !reg_error;

  assign dout_7_re = addr_hit[57] & reg_re & !reg_error;

  assign dout_8_re = addr_hit[58] & reg_re & !reg_error;

  assign dout_9_re = addr_hit[59] & reg_re & !reg_error;

  assign dout_10_re = addr_hit[60] & reg_re & !reg_error;

  assign dout_11_re = addr_hit[61] & reg_re & !reg_error;

  assign dout_12_re = addr_hit[62] & reg_re & !reg_error;

  assign dout_13_re = addr_hit[63] & reg_re & !reg_error;

  assign dout_14_re = addr_hit[64] & reg_re & !reg_error;

  assign dout_15_re = addr_hit[65] & reg_re & !reg_error;

  assign dout_16_re = addr_hit[66] & reg_re & !reg_error;

  assign dout_17_re = addr_hit[67] & reg_re & !reg_error;

  assign dout_18_re = addr_hit[68] & reg_re & !reg_error;

  assign dout_19_re = addr_hit[69] & reg_re & !reg_error;

  assign dout_20_re = addr_hit[70] & reg_re & !reg_error;

  assign dout_21_re = addr_hit[71] & reg_re & !reg_error;

  assign dout_22_re = addr_hit[72] & reg_re & !reg_error;

  assign dout_23_re = addr_hit[73] & reg_re & !reg_error;

  assign dout_24_re = addr_hit[74] & reg_re & !reg_error;

  assign dout_25_re = addr_hit[75] & reg_re & !reg_error;

  assign dout_26_re = addr_hit[76] & reg_re & !reg_error;

  assign dout_27_re = addr_hit[77] & reg_re & !reg_error;

  assign dout_28_re = addr_hit[78] & reg_re & !reg_error;

  assign dout_29_re = addr_hit[79] & reg_re & !reg_error;

  assign dout_30_re = addr_hit[80] & reg_re & !reg_error;

  assign dout_31_re = addr_hit[81] & reg_re & !reg_error;

  assign dout_32_re = addr_hit[82] & reg_re & !reg_error;

  assign dout_33_re = addr_hit[83] & reg_re & !reg_error;

  assign dout_34_re = addr_hit[84] & reg_re & !reg_error;

  assign dout_35_re = addr_hit[85] & reg_re & !reg_error;

  assign dout_36_re = addr_hit[86] & reg_re & !reg_error;

  assign dout_37_re = addr_hit[87] & reg_re & !reg_error;

  assign dout_38_re = addr_hit[88] & reg_re & !reg_error;

  assign dout_39_re = addr_hit[89] & reg_re & !reg_error;

  assign dout_40_re = addr_hit[90] & reg_re & !reg_error;

  assign dout_41_re = addr_hit[91] & reg_re & !reg_error;

  assign dout_42_re = addr_hit[92] & reg_re & !reg_error;

  assign dout_43_re = addr_hit[93] & reg_re & !reg_error;

  assign dout_44_re = addr_hit[94] & reg_re & !reg_error;

  assign dout_45_re = addr_hit[95] & reg_re & !reg_error;

  assign dout_46_re = addr_hit[96] & reg_re & !reg_error;

  assign dout_47_re = addr_hit[97] & reg_re & !reg_error;

  assign dout_48_re = addr_hit[98] & reg_re & !reg_error;

  assign dout_49_re = addr_hit[99] & reg_re & !reg_error;

  // Read data return
  always_comb begin
    reg_rdata_next = '0;
    unique case (1'b1)
      addr_hit[0]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[1]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[2]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[3]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[4]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[5]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[6]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[7]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[8]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[9]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[10]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[11]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[12]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[13]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[14]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[15]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[16]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[17]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[18]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[19]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[20]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[21]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[22]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[23]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[24]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[25]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[26]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[27]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[28]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[29]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[30]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[31]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[32]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[33]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[34]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[35]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[36]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[37]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[38]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[39]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[40]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[41]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[42]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[43]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[44]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[45]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[46]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[47]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[48]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[49]: begin
        reg_rdata_next[31:0] = '0;
      end

      addr_hit[50]: begin
        reg_rdata_next[31:0] = dout_0_qs;
      end

      addr_hit[51]: begin
        reg_rdata_next[31:0] = dout_1_qs;
      end

      addr_hit[52]: begin
        reg_rdata_next[31:0] = dout_2_qs;
      end

      addr_hit[53]: begin
        reg_rdata_next[31:0] = dout_3_qs;
      end

      addr_hit[54]: begin
        reg_rdata_next[31:0] = dout_4_qs;
      end

      addr_hit[55]: begin
        reg_rdata_next[31:0] = dout_5_qs;
      end

      addr_hit[56]: begin
        reg_rdata_next[31:0] = dout_6_qs;
      end

      addr_hit[57]: begin
        reg_rdata_next[31:0] = dout_7_qs;
      end

      addr_hit[58]: begin
        reg_rdata_next[31:0] = dout_8_qs;
      end

      addr_hit[59]: begin
        reg_rdata_next[31:0] = dout_9_qs;
      end

      addr_hit[60]: begin
        reg_rdata_next[31:0] = dout_10_qs;
      end

      addr_hit[61]: begin
        reg_rdata_next[31:0] = dout_11_qs;
      end

      addr_hit[62]: begin
        reg_rdata_next[31:0] = dout_12_qs;
      end

      addr_hit[63]: begin
        reg_rdata_next[31:0] = dout_13_qs;
      end

      addr_hit[64]: begin
        reg_rdata_next[31:0] = dout_14_qs;
      end

      addr_hit[65]: begin
        reg_rdata_next[31:0] = dout_15_qs;
      end

      addr_hit[66]: begin
        reg_rdata_next[31:0] = dout_16_qs;
      end

      addr_hit[67]: begin
        reg_rdata_next[31:0] = dout_17_qs;
      end

      addr_hit[68]: begin
        reg_rdata_next[31:0] = dout_18_qs;
      end

      addr_hit[69]: begin
        reg_rdata_next[31:0] = dout_19_qs;
      end

      addr_hit[70]: begin
        reg_rdata_next[31:0] = dout_20_qs;
      end

      addr_hit[71]: begin
        reg_rdata_next[31:0] = dout_21_qs;
      end

      addr_hit[72]: begin
        reg_rdata_next[31:0] = dout_22_qs;
      end

      addr_hit[73]: begin
        reg_rdata_next[31:0] = dout_23_qs;
      end

      addr_hit[74]: begin
        reg_rdata_next[31:0] = dout_24_qs;
      end

      addr_hit[75]: begin
        reg_rdata_next[31:0] = dout_25_qs;
      end

      addr_hit[76]: begin
        reg_rdata_next[31:0] = dout_26_qs;
      end

      addr_hit[77]: begin
        reg_rdata_next[31:0] = dout_27_qs;
      end

      addr_hit[78]: begin
        reg_rdata_next[31:0] = dout_28_qs;
      end

      addr_hit[79]: begin
        reg_rdata_next[31:0] = dout_29_qs;
      end

      addr_hit[80]: begin
        reg_rdata_next[31:0] = dout_30_qs;
      end

      addr_hit[81]: begin
        reg_rdata_next[31:0] = dout_31_qs;
      end

      addr_hit[82]: begin
        reg_rdata_next[31:0] = dout_32_qs;
      end

      addr_hit[83]: begin
        reg_rdata_next[31:0] = dout_33_qs;
      end

      addr_hit[84]: begin
        reg_rdata_next[31:0] = dout_34_qs;
      end

      addr_hit[85]: begin
        reg_rdata_next[31:0] = dout_35_qs;
      end

      addr_hit[86]: begin
        reg_rdata_next[31:0] = dout_36_qs;
      end

      addr_hit[87]: begin
        reg_rdata_next[31:0] = dout_37_qs;
      end

      addr_hit[88]: begin
        reg_rdata_next[31:0] = dout_38_qs;
      end

      addr_hit[89]: begin
        reg_rdata_next[31:0] = dout_39_qs;
      end

      addr_hit[90]: begin
        reg_rdata_next[31:0] = dout_40_qs;
      end

      addr_hit[91]: begin
        reg_rdata_next[31:0] = dout_41_qs;
      end

      addr_hit[92]: begin
        reg_rdata_next[31:0] = dout_42_qs;
      end

      addr_hit[93]: begin
        reg_rdata_next[31:0] = dout_43_qs;
      end

      addr_hit[94]: begin
        reg_rdata_next[31:0] = dout_44_qs;
      end

      addr_hit[95]: begin
        reg_rdata_next[31:0] = dout_45_qs;
      end

      addr_hit[96]: begin
        reg_rdata_next[31:0] = dout_46_qs;
      end

      addr_hit[97]: begin
        reg_rdata_next[31:0] = dout_47_qs;
      end

      addr_hit[98]: begin
        reg_rdata_next[31:0] = dout_48_qs;
      end

      addr_hit[99]: begin
        reg_rdata_next[31:0] = dout_49_qs;
      end

      default: begin
        reg_rdata_next = '1;
      end
    endcase
  end

  // Unused signal tieoff

  // wdata / byte enable are not always fully used
  // add a blanket unused statement to handle lint waivers
  logic unused_wdata;
  logic unused_be;
  assign unused_wdata = ^reg_wdata;
  assign unused_be = ^reg_be;

  // Assertions for Register Interface
  `ASSERT(en2addrHit, (reg_we || reg_re) |-> $onehot0(addr_hit))

endmodule

module keccak_data_reg_top_intf
#(
  parameter int AW = 9,
  localparam int DW = 32
) (
  input logic clk_i,
  input logic rst_ni,
  REG_BUS.in  regbus_slave,
  // To HW
  output keccak_data_reg_pkg::keccak_data_reg2hw_t reg2hw, // Write
  input  keccak_data_reg_pkg::keccak_data_hw2reg_t hw2reg, // Read
  // Config
  input devmode_i // If 1, explicit error return for unmapped register access
);
 localparam int unsigned STRB_WIDTH = DW/8;

`include "register_interface/typedef.svh"
`include "register_interface/assign.svh"

  // Define structs for reg_bus
  typedef logic [AW-1:0] addr_t;
  typedef logic [DW-1:0] data_t;
  typedef logic [STRB_WIDTH-1:0] strb_t;
  `REG_BUS_TYPEDEF_ALL(reg_bus, addr_t, data_t, strb_t)

  reg_bus_req_t s_reg_req;
  reg_bus_rsp_t s_reg_rsp;
  
  // Assign SV interface to structs
  `REG_BUS_ASSIGN_TO_REQ(s_reg_req, regbus_slave)
  `REG_BUS_ASSIGN_FROM_RSP(regbus_slave, s_reg_rsp)

  

  keccak_data_reg_top #(
    .reg_req_t(reg_bus_req_t),
    .reg_rsp_t(reg_bus_rsp_t),
    .AW(AW)
  ) i_regs (
    .clk_i,
    .rst_ni,
    .reg_req_i(s_reg_req),
    .reg_rsp_o(s_reg_rsp),
    .reg2hw, // Write
    .hw2reg, // Read
    .devmode_i
  );
  
endmodule


