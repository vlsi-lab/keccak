//////////////////////////////////////////////////////////////////////////////////////////
// Authors:      Alessandra Dolmeta - alessandra.dolmeta@polito.it                      //
//               Valeria Piscopo    - valeria.piscopo@polito.it                         //
//               Mattia Mirigaldi    - mattia.mirigaldi@polito.it                       //
// Language:     SystemVerilog                                                          //
// Based on the designed of Michal Peeters and Gilles Van Assche.                       //
//                                                                                      //
//////////////////////////////////////////////////////////////////////////////////////////

// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package keccak_ctrl_reg_pkg;

  // Address widths within the block
  parameter int BlockAw = 3;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    logic        q;
  } keccak_ctrl_reg2hw_ctrl_reg_t;

  typedef struct packed {
    logic        d;
    logic        de;
  } keccak_ctrl_hw2reg_status_reg_t;

  // Register -> HW type
  typedef struct packed {
    keccak_ctrl_reg2hw_ctrl_reg_t ctrl; // [0:0]
  } keccak_ctrl_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    keccak_ctrl_hw2reg_status_reg_t status; // [1:0]
  } keccak_ctrl_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] KECCAK_CTRL_CTRL_OFFSET = 3'h 0;
  parameter logic [BlockAw-1:0] KECCAK_CTRL_STATUS_OFFSET = 3'h 4;

  // Register index
  typedef enum int {
    KECCAK_CTRL_CTRL,
    KECCAK_CTRL_STATUS
  } keccak_ctrl_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] KECCAK_CTRL_PERMIT [2] = '{
    4'b 0001, // index[0] KECCAK_CTRL_CTRL
    4'b 0001  // index[1] KECCAK_CTRL_STATUS
  };

endpackage

