//////////////////////////////////////////////////////////////////////////////////////////
// Authors:      Alessandra Dolmeta - alessandra.dolmeta@polito.it                      //
//               Valeria Piscopo    - valeria.piscopo@polito.it                         //
//               Mattia Mirigaldi    - mattia.mirigaldi@polito.it                       //
// Language:     SystemVerilog                                                          //
// Based on the designed of Michal Peeters and Gilles Van Assche.                       //
//                                                                                      //
//////////////////////////////////////////////////////////////////////////////////////////

// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// Register Package auto-generated by `reggen` containing data structure

package keccak_data_reg_pkg;

  // Address widths within the block
  parameter int BlockAw = 9;

  ////////////////////////////
  // Typedefs for registers //
  ////////////////////////////

  typedef struct packed {
    logic [31:0] q;
  } keccak_data_reg2hw_din_mreg_t;

  typedef struct packed {
    logic [31:0] d;
  } keccak_data_hw2reg_dout_mreg_t;

  // Register -> HW type
  typedef struct packed {
    keccak_data_reg2hw_din_mreg_t [49:0] din; // [1599:0]
  } keccak_data_reg2hw_t;

  // HW -> register type
  typedef struct packed {
    keccak_data_hw2reg_dout_mreg_t [49:0] dout; // [1599:0]
  } keccak_data_hw2reg_t;

  // Register offsets
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_0_OFFSET = 9'h 0;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_1_OFFSET = 9'h 4;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_2_OFFSET = 9'h 8;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_3_OFFSET = 9'h c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_4_OFFSET = 9'h 10;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_5_OFFSET = 9'h 14;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_6_OFFSET = 9'h 18;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_7_OFFSET = 9'h 1c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_8_OFFSET = 9'h 20;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_9_OFFSET = 9'h 24;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_10_OFFSET = 9'h 28;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_11_OFFSET = 9'h 2c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_12_OFFSET = 9'h 30;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_13_OFFSET = 9'h 34;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_14_OFFSET = 9'h 38;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_15_OFFSET = 9'h 3c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_16_OFFSET = 9'h 40;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_17_OFFSET = 9'h 44;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_18_OFFSET = 9'h 48;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_19_OFFSET = 9'h 4c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_20_OFFSET = 9'h 50;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_21_OFFSET = 9'h 54;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_22_OFFSET = 9'h 58;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_23_OFFSET = 9'h 5c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_24_OFFSET = 9'h 60;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_25_OFFSET = 9'h 64;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_26_OFFSET = 9'h 68;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_27_OFFSET = 9'h 6c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_28_OFFSET = 9'h 70;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_29_OFFSET = 9'h 74;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_30_OFFSET = 9'h 78;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_31_OFFSET = 9'h 7c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_32_OFFSET = 9'h 80;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_33_OFFSET = 9'h 84;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_34_OFFSET = 9'h 88;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_35_OFFSET = 9'h 8c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_36_OFFSET = 9'h 90;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_37_OFFSET = 9'h 94;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_38_OFFSET = 9'h 98;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_39_OFFSET = 9'h 9c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_40_OFFSET = 9'h a0;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_41_OFFSET = 9'h a4;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_42_OFFSET = 9'h a8;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_43_OFFSET = 9'h ac;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_44_OFFSET = 9'h b0;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_45_OFFSET = 9'h b4;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_46_OFFSET = 9'h b8;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_47_OFFSET = 9'h bc;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_48_OFFSET = 9'h c0;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DIN_49_OFFSET = 9'h c4;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_0_OFFSET = 9'h c8;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_1_OFFSET = 9'h cc;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_2_OFFSET = 9'h d0;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_3_OFFSET = 9'h d4;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_4_OFFSET = 9'h d8;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_5_OFFSET = 9'h dc;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_6_OFFSET = 9'h e0;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_7_OFFSET = 9'h e4;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_8_OFFSET = 9'h e8;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_9_OFFSET = 9'h ec;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_10_OFFSET = 9'h f0;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_11_OFFSET = 9'h f4;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_12_OFFSET = 9'h f8;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_13_OFFSET = 9'h fc;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_14_OFFSET = 9'h 100;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_15_OFFSET = 9'h 104;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_16_OFFSET = 9'h 108;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_17_OFFSET = 9'h 10c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_18_OFFSET = 9'h 110;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_19_OFFSET = 9'h 114;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_20_OFFSET = 9'h 118;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_21_OFFSET = 9'h 11c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_22_OFFSET = 9'h 120;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_23_OFFSET = 9'h 124;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_24_OFFSET = 9'h 128;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_25_OFFSET = 9'h 12c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_26_OFFSET = 9'h 130;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_27_OFFSET = 9'h 134;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_28_OFFSET = 9'h 138;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_29_OFFSET = 9'h 13c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_30_OFFSET = 9'h 140;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_31_OFFSET = 9'h 144;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_32_OFFSET = 9'h 148;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_33_OFFSET = 9'h 14c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_34_OFFSET = 9'h 150;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_35_OFFSET = 9'h 154;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_36_OFFSET = 9'h 158;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_37_OFFSET = 9'h 15c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_38_OFFSET = 9'h 160;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_39_OFFSET = 9'h 164;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_40_OFFSET = 9'h 168;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_41_OFFSET = 9'h 16c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_42_OFFSET = 9'h 170;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_43_OFFSET = 9'h 174;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_44_OFFSET = 9'h 178;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_45_OFFSET = 9'h 17c;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_46_OFFSET = 9'h 180;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_47_OFFSET = 9'h 184;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_48_OFFSET = 9'h 188;
  parameter logic [BlockAw-1:0] KECCAK_DATA_DOUT_49_OFFSET = 9'h 18c;

  // Reset values for hwext registers and their fields
  parameter logic [31:0] KECCAK_DATA_DOUT_0_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_1_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_2_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_3_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_4_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_5_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_6_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_7_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_8_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_9_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_10_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_11_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_12_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_13_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_14_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_15_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_16_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_17_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_18_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_19_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_20_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_21_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_22_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_23_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_24_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_25_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_26_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_27_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_28_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_29_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_30_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_31_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_32_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_33_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_34_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_35_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_36_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_37_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_38_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_39_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_40_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_41_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_42_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_43_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_44_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_45_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_46_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_47_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_48_RESVAL = 32'h 0;
  parameter logic [31:0] KECCAK_DATA_DOUT_49_RESVAL = 32'h 0;

  // Register index
  typedef enum int {
    KECCAK_DATA_DIN_0,
    KECCAK_DATA_DIN_1,
    KECCAK_DATA_DIN_2,
    KECCAK_DATA_DIN_3,
    KECCAK_DATA_DIN_4,
    KECCAK_DATA_DIN_5,
    KECCAK_DATA_DIN_6,
    KECCAK_DATA_DIN_7,
    KECCAK_DATA_DIN_8,
    KECCAK_DATA_DIN_9,
    KECCAK_DATA_DIN_10,
    KECCAK_DATA_DIN_11,
    KECCAK_DATA_DIN_12,
    KECCAK_DATA_DIN_13,
    KECCAK_DATA_DIN_14,
    KECCAK_DATA_DIN_15,
    KECCAK_DATA_DIN_16,
    KECCAK_DATA_DIN_17,
    KECCAK_DATA_DIN_18,
    KECCAK_DATA_DIN_19,
    KECCAK_DATA_DIN_20,
    KECCAK_DATA_DIN_21,
    KECCAK_DATA_DIN_22,
    KECCAK_DATA_DIN_23,
    KECCAK_DATA_DIN_24,
    KECCAK_DATA_DIN_25,
    KECCAK_DATA_DIN_26,
    KECCAK_DATA_DIN_27,
    KECCAK_DATA_DIN_28,
    KECCAK_DATA_DIN_29,
    KECCAK_DATA_DIN_30,
    KECCAK_DATA_DIN_31,
    KECCAK_DATA_DIN_32,
    KECCAK_DATA_DIN_33,
    KECCAK_DATA_DIN_34,
    KECCAK_DATA_DIN_35,
    KECCAK_DATA_DIN_36,
    KECCAK_DATA_DIN_37,
    KECCAK_DATA_DIN_38,
    KECCAK_DATA_DIN_39,
    KECCAK_DATA_DIN_40,
    KECCAK_DATA_DIN_41,
    KECCAK_DATA_DIN_42,
    KECCAK_DATA_DIN_43,
    KECCAK_DATA_DIN_44,
    KECCAK_DATA_DIN_45,
    KECCAK_DATA_DIN_46,
    KECCAK_DATA_DIN_47,
    KECCAK_DATA_DIN_48,
    KECCAK_DATA_DIN_49,
    KECCAK_DATA_DOUT_0,
    KECCAK_DATA_DOUT_1,
    KECCAK_DATA_DOUT_2,
    KECCAK_DATA_DOUT_3,
    KECCAK_DATA_DOUT_4,
    KECCAK_DATA_DOUT_5,
    KECCAK_DATA_DOUT_6,
    KECCAK_DATA_DOUT_7,
    KECCAK_DATA_DOUT_8,
    KECCAK_DATA_DOUT_9,
    KECCAK_DATA_DOUT_10,
    KECCAK_DATA_DOUT_11,
    KECCAK_DATA_DOUT_12,
    KECCAK_DATA_DOUT_13,
    KECCAK_DATA_DOUT_14,
    KECCAK_DATA_DOUT_15,
    KECCAK_DATA_DOUT_16,
    KECCAK_DATA_DOUT_17,
    KECCAK_DATA_DOUT_18,
    KECCAK_DATA_DOUT_19,
    KECCAK_DATA_DOUT_20,
    KECCAK_DATA_DOUT_21,
    KECCAK_DATA_DOUT_22,
    KECCAK_DATA_DOUT_23,
    KECCAK_DATA_DOUT_24,
    KECCAK_DATA_DOUT_25,
    KECCAK_DATA_DOUT_26,
    KECCAK_DATA_DOUT_27,
    KECCAK_DATA_DOUT_28,
    KECCAK_DATA_DOUT_29,
    KECCAK_DATA_DOUT_30,
    KECCAK_DATA_DOUT_31,
    KECCAK_DATA_DOUT_32,
    KECCAK_DATA_DOUT_33,
    KECCAK_DATA_DOUT_34,
    KECCAK_DATA_DOUT_35,
    KECCAK_DATA_DOUT_36,
    KECCAK_DATA_DOUT_37,
    KECCAK_DATA_DOUT_38,
    KECCAK_DATA_DOUT_39,
    KECCAK_DATA_DOUT_40,
    KECCAK_DATA_DOUT_41,
    KECCAK_DATA_DOUT_42,
    KECCAK_DATA_DOUT_43,
    KECCAK_DATA_DOUT_44,
    KECCAK_DATA_DOUT_45,
    KECCAK_DATA_DOUT_46,
    KECCAK_DATA_DOUT_47,
    KECCAK_DATA_DOUT_48,
    KECCAK_DATA_DOUT_49
  } keccak_data_id_e;

  // Register width information to check illegal writes
  parameter logic [3:0] KECCAK_DATA_PERMIT [100] = '{
    4'b 1111, // index[ 0] KECCAK_DATA_DIN_0
    4'b 1111, // index[ 1] KECCAK_DATA_DIN_1
    4'b 1111, // index[ 2] KECCAK_DATA_DIN_2
    4'b 1111, // index[ 3] KECCAK_DATA_DIN_3
    4'b 1111, // index[ 4] KECCAK_DATA_DIN_4
    4'b 1111, // index[ 5] KECCAK_DATA_DIN_5
    4'b 1111, // index[ 6] KECCAK_DATA_DIN_6
    4'b 1111, // index[ 7] KECCAK_DATA_DIN_7
    4'b 1111, // index[ 8] KECCAK_DATA_DIN_8
    4'b 1111, // index[ 9] KECCAK_DATA_DIN_9
    4'b 1111, // index[10] KECCAK_DATA_DIN_10
    4'b 1111, // index[11] KECCAK_DATA_DIN_11
    4'b 1111, // index[12] KECCAK_DATA_DIN_12
    4'b 1111, // index[13] KECCAK_DATA_DIN_13
    4'b 1111, // index[14] KECCAK_DATA_DIN_14
    4'b 1111, // index[15] KECCAK_DATA_DIN_15
    4'b 1111, // index[16] KECCAK_DATA_DIN_16
    4'b 1111, // index[17] KECCAK_DATA_DIN_17
    4'b 1111, // index[18] KECCAK_DATA_DIN_18
    4'b 1111, // index[19] KECCAK_DATA_DIN_19
    4'b 1111, // index[20] KECCAK_DATA_DIN_20
    4'b 1111, // index[21] KECCAK_DATA_DIN_21
    4'b 1111, // index[22] KECCAK_DATA_DIN_22
    4'b 1111, // index[23] KECCAK_DATA_DIN_23
    4'b 1111, // index[24] KECCAK_DATA_DIN_24
    4'b 1111, // index[25] KECCAK_DATA_DIN_25
    4'b 1111, // index[26] KECCAK_DATA_DIN_26
    4'b 1111, // index[27] KECCAK_DATA_DIN_27
    4'b 1111, // index[28] KECCAK_DATA_DIN_28
    4'b 1111, // index[29] KECCAK_DATA_DIN_29
    4'b 1111, // index[30] KECCAK_DATA_DIN_30
    4'b 1111, // index[31] KECCAK_DATA_DIN_31
    4'b 1111, // index[32] KECCAK_DATA_DIN_32
    4'b 1111, // index[33] KECCAK_DATA_DIN_33
    4'b 1111, // index[34] KECCAK_DATA_DIN_34
    4'b 1111, // index[35] KECCAK_DATA_DIN_35
    4'b 1111, // index[36] KECCAK_DATA_DIN_36
    4'b 1111, // index[37] KECCAK_DATA_DIN_37
    4'b 1111, // index[38] KECCAK_DATA_DIN_38
    4'b 1111, // index[39] KECCAK_DATA_DIN_39
    4'b 1111, // index[40] KECCAK_DATA_DIN_40
    4'b 1111, // index[41] KECCAK_DATA_DIN_41
    4'b 1111, // index[42] KECCAK_DATA_DIN_42
    4'b 1111, // index[43] KECCAK_DATA_DIN_43
    4'b 1111, // index[44] KECCAK_DATA_DIN_44
    4'b 1111, // index[45] KECCAK_DATA_DIN_45
    4'b 1111, // index[46] KECCAK_DATA_DIN_46
    4'b 1111, // index[47] KECCAK_DATA_DIN_47
    4'b 1111, // index[48] KECCAK_DATA_DIN_48
    4'b 1111, // index[49] KECCAK_DATA_DIN_49
    4'b 1111, // index[50] KECCAK_DATA_DOUT_0
    4'b 1111, // index[51] KECCAK_DATA_DOUT_1
    4'b 1111, // index[52] KECCAK_DATA_DOUT_2
    4'b 1111, // index[53] KECCAK_DATA_DOUT_3
    4'b 1111, // index[54] KECCAK_DATA_DOUT_4
    4'b 1111, // index[55] KECCAK_DATA_DOUT_5
    4'b 1111, // index[56] KECCAK_DATA_DOUT_6
    4'b 1111, // index[57] KECCAK_DATA_DOUT_7
    4'b 1111, // index[58] KECCAK_DATA_DOUT_8
    4'b 1111, // index[59] KECCAK_DATA_DOUT_9
    4'b 1111, // index[60] KECCAK_DATA_DOUT_10
    4'b 1111, // index[61] KECCAK_DATA_DOUT_11
    4'b 1111, // index[62] KECCAK_DATA_DOUT_12
    4'b 1111, // index[63] KECCAK_DATA_DOUT_13
    4'b 1111, // index[64] KECCAK_DATA_DOUT_14
    4'b 1111, // index[65] KECCAK_DATA_DOUT_15
    4'b 1111, // index[66] KECCAK_DATA_DOUT_16
    4'b 1111, // index[67] KECCAK_DATA_DOUT_17
    4'b 1111, // index[68] KECCAK_DATA_DOUT_18
    4'b 1111, // index[69] KECCAK_DATA_DOUT_19
    4'b 1111, // index[70] KECCAK_DATA_DOUT_20
    4'b 1111, // index[71] KECCAK_DATA_DOUT_21
    4'b 1111, // index[72] KECCAK_DATA_DOUT_22
    4'b 1111, // index[73] KECCAK_DATA_DOUT_23
    4'b 1111, // index[74] KECCAK_DATA_DOUT_24
    4'b 1111, // index[75] KECCAK_DATA_DOUT_25
    4'b 1111, // index[76] KECCAK_DATA_DOUT_26
    4'b 1111, // index[77] KECCAK_DATA_DOUT_27
    4'b 1111, // index[78] KECCAK_DATA_DOUT_28
    4'b 1111, // index[79] KECCAK_DATA_DOUT_29
    4'b 1111, // index[80] KECCAK_DATA_DOUT_30
    4'b 1111, // index[81] KECCAK_DATA_DOUT_31
    4'b 1111, // index[82] KECCAK_DATA_DOUT_32
    4'b 1111, // index[83] KECCAK_DATA_DOUT_33
    4'b 1111, // index[84] KECCAK_DATA_DOUT_34
    4'b 1111, // index[85] KECCAK_DATA_DOUT_35
    4'b 1111, // index[86] KECCAK_DATA_DOUT_36
    4'b 1111, // index[87] KECCAK_DATA_DOUT_37
    4'b 1111, // index[88] KECCAK_DATA_DOUT_38
    4'b 1111, // index[89] KECCAK_DATA_DOUT_39
    4'b 1111, // index[90] KECCAK_DATA_DOUT_40
    4'b 1111, // index[91] KECCAK_DATA_DOUT_41
    4'b 1111, // index[92] KECCAK_DATA_DOUT_42
    4'b 1111, // index[93] KECCAK_DATA_DOUT_43
    4'b 1111, // index[94] KECCAK_DATA_DOUT_44
    4'b 1111, // index[95] KECCAK_DATA_DOUT_45
    4'b 1111, // index[96] KECCAK_DATA_DOUT_46
    4'b 1111, // index[97] KECCAK_DATA_DOUT_47
    4'b 1111, // index[98] KECCAK_DATA_DOUT_48
    4'b 1111  // index[99] KECCAK_DATA_DOUT_49
  };

endpackage

